Vim�UnDo� ���r��u�����ݴ@a3����	ǉ��d   8   $        $display("rsort =  %p",res);   0   "                   aL    _�                             ����                                                                                                                                                                                                                                                                                                                                                            aE{�     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aE{�     �                     int array[9]='{};5�_�                       /    ����                                                                                                                                                                                                                                                                                                                                                            aE{�     �                 /    int array[9]='{12,14,32,45,56,76,47,72,94};5�_�                            ����                                                                                                                                                                                                                                                                                                                                                            aE{�     �                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aE|     �                       res = array.find()5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aE|     �                       res = array.find(x)5�_�                       "    ����                                                                                                                                                                                                                                                                                                                                                            aE|     �               #        res = array.find(x) with ()5�_�      	                 &    ����                                                                                                                                                                                                                                                                                                                                                            aE|     �      	         &        res = array.find(x) with (x>3)5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                            aE|     �      	   	              $display()5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                            aE|     �      	   	              $display();5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                            aE|     �      	   	              $display("");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aE|     �      	   	              $display("find()");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aE|!     �      	   	              $display("find(x)");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aE|&     �      	   	      !        $display("find(x) : %p");5�_�                       %    ����                                                                                                                                                                                                                                                                                                                                                            aE|)     �         	      %        $display("find(x) : %p",res);5�_�                    
        ����                                                                                                                                                                                                                                                                                                                                                            aE|7     �   	             �   
          5�_�                    
        ����                                                                                                                                                                                                                                                                                                                                                            aE|8     �   	             �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                            aE|8     �   	              �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                            aE|9     �   	               �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                            aE|:     �   	                �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                            aE|:     �   	                 �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                            aE|:     �   	                  �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                            aE|;     �   	                   �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                            aE|<     �   	                    �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                            aE|@     �   	            	         �   
          5�_�                    
   	    ����                                                                                                                                                                                                                                                                                                                                                            aE|@     �   	            
          �   
          5�_�                    
   
    ����                                                                                                                                                                                                                                                                                                                                                            aE|A     �   	                       �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                     	           v       aE|p     �   	                        �   
          5�_�                           ����                                                                                                                                                                                                                                                                                                                                     	           v       aE|s     �                    �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                     	           v       aE|z     �                �             5�_�                             ����                                                                                                                                                                                                                                                                                                                                     	           v       aE||     �                �             5�_�      !                       ����                                                                                                                                                                                                                                                                                                                                     	           v       aE|�     �                �             5�_�       "           !   
       ����                                                                                                                                                                                                                                                                                                                                     	           v       aE|�    �   	            (         res = array.find(x) with (x>3);5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                            aE��     �               !  res = array.find(x) with (x>3);5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                            aE��     �               !  res = array.find(x) with (x>3);5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                            aE��     �               !  res = array.find(x) with (x>3);5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                            aE��     �               &       res = array.find(x) with (x>3);5�_�   %   (           &   
   '    ����                                                                                                                                                                                                                                                                                                                                                            aE��     �   	            '        res = array.find(x) with (x>3);5�_�   &   )   '       (           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                 '        res = array.find(x) with (x>3);   %        $display("find(x) : %p",res);       '        res = array.find(x) with (x>3);   %        $display("find(x) : %p",res);       '        res = array.find(x) with (x>3);   %        $display("find(x) : %p",res);       '        res = array.find(x) with (x>3);   %        $display("find(x) : %p",res);       '        res = array.find(x) with (x>3);   %        $display("find(x) : %p",res);       '        res = array.find(x) with (x>3);   %        $display("find(x) : %p",res);               end5�_�   (   *           )           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                     end5�_�   )   +           *           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                       res=array.find()5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                       res=array.find(x)5�_�   ,   .           -           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �               !        res=array.find(x) with ()5�_�   -   /           .      $    ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �      	         $        res=array.find(x) with (x>3)5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �      	   	              $display()5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �      	   	              $display("")5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�      �      	   	              $display("");5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�     �      	   	              $display("finc()");5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�     �      	   	              $display("finc(x)");5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�     �      	   	      !        $display("finc(x) : %p");5�_�   4   6           5      %    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�     �         	      %        $display("finc(x) : %p",res);5�_�   5   7           6   
        ����                                                                                                                                                                                                                                                                                                                                     
           v       aE�     �   	             �   
          5�_�   6   8           7   
        ����                                                                                                                                                                                                                                                                                                                                     
           v       aE�     �   	             res=array.find(x) with (x>3);5�_�   7   9           8   
   	    ����                                                                                                                                                                                                                                                                                                                                     
           v       aE�    �   	            &         res=array.find(x) with (x>3);5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                            aE�7     �                     end5�_�   9   ;           :   
       ����                                                                                                                                                                                                                                                                                                                                                            aE�S     �   	            %        res=array.find(x) with (x>3);5�_�   :   <           ;   
       ����                                                                                                                                                                                                                                                                                                                                                            aE�U     �   	            #        res=array.find) with (x>3);5�_�   ;   =           <   
   &    ����                                                                                                                                                                                                                                                                                                                                                            aE�]     �   	            (        res=array.find_index with (x>3);5�_�   <   >           =   
   *    ����                                                                                                                                                                                                                                                                                                                                                            aE�b     �   	            -        res=array.find_index with (item ==4);5�_�   =   ?           >   
   ,    ����                                                                                                                                                                                                                                                                                                                                                            aE�d     �   	            .        res=array.find_index with (item == 4);5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                            aE�l     �      	         %        $display("finc(x) : %p",res);5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                            aE�r     �   
            %        $display("finc(x) : %p",res);5�_�   @   B           A      #    ����                                                                                                                                                                                                                                                                                                                                                            aE�|     �   
            %        $display("find(x) : %p",res);5�_�   A   C           B          ����                                                                                                                                                                                                                                                                                                                                                            aE��     �   
            -        $display("find(x) : %p",res[%0d]=32);5�_�   B   D           C          ����                                                                                                                                                                                                                                                                                                                                                            aE��     �   
            *        $display("find(x) : ,res[%0d]=32);5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                                                            aE��     �   
            )        $display("find(x) : res[%0d]=32);5�_�   D   F           E      *    ����                                                                                                                                                                                                                                                                                                                                                            aE��     �   
            ,        $display("find_index : res[%0d]=32);5�_�   E   G           F      3    ����                                                                                                                                                                                                                                                                                                                                                            aE��     �   
            3        $display("find_index : res[%0d]=32,res[0]);5�_�   F   H           G           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                       �             5�_�   H   J           I      	    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �               0         res=array.find_index with (item == 32);5�_�   I   K           J           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                       �             5�_�   K   M           L      	    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �               0         res=array.find_index with (item == 32);5�_�   L   N           M           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                       �             5�_�   N   P           O      	    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �               0         res=array.find_index with (item == 32);5�_�   O   Q           P           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                5�_�   P   R           Q           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                    �                    �                    �                    �                    �                    �                5�_�   Q   S           R           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                5�_�   R   T           S           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                �             5�_�   S   U           T           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �               ( res=array.find_index with (item == 32);5�_�   T   V           U      	    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �               0         res=array.find_index with (item == 32);5�_�   U   W           V           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                5�_�   V   X           W           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                5�_�   W   Y           X           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                5�_�   X   Z           Y           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                5�_�   Y   [           Z           ����                                                                                                                                                                                                                                                                                                                           
                     v       aE��     �                    �                    �                    �                5�_�   Z   \           [      *    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�     �   
            3        $display("find_index : res[%0d]=32,res[0]);5�_�   [   ]           \          ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�     �               /        res=array.find_index with (item == 32);5�_�   \   ^           ]      *    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�!     �               /        res=array.find_first with (item == 32);5�_�   ]   _           ^      8    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�/     �               :        res=array.find_first with (item <15 & item >= 32);5�_�   ^   `           _      5    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�>     �               8        res=array.find_first with (item <15 & item >= );5�_�   _   a           `      8    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�D     �               :        res=array.find_first with (item <15 & item >=13 );5�_�   `   b           a          ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�M     �               3        $display("find_index : res[%0d]=32,res[0]);5�_�   a   c           b      *    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�b     �               3        $display("find_first : res[%0d]=32,res[0]);5�_�   b   d           c      *    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�c     �               4        $display("find_first : res[%0d]=32",res[0]);5�_�   c   e           d      )    ����                                                                                                                                                                                                                                                                                                                           
                     v       aE�m     �               +        $display("find_first : %p",res[0]);5�_�   d   f           e           ����                                                                                                                                                                                                                                                                                                                                         %       v   %    aE�u     �            	       /        res=array.find_index with (item == 32);   3        $display("find_index : res[%0d]=32,res[0]);       /        res=array.find_index with (item == 32);   3        $display("find_index : res[%0d]=32,res[0]);       /        res=array.find_index with (item == 32);   3        $display("find_index : res[%0d]=32,res[0]);5�_�   e   g           f           ����                                                                                                                                                                                                                                                                                                                                                 v        aE�x     �               ]=32,res[0]);           end5�_�   f   h           g           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                   end5�_�   g   i           h           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                5�_�   h   j           i           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                5�_�   i   k           j          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                       5�_�   j   l           k          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �               	         �             5�_�   k   m           l           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                 5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                 5�_�   m   o           n          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �               	         5�_�   n   p           o          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �             �             5�_�   o   q           p           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �             �             5�_�   p   s           q           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �               
          �             5�_�   q   t   r       s           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �               
          �             5�_�   s   u           t           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                 5�_�   t   v           u          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                	         5�_�   u   w           v           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                 5�_�   v   x           w          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                	         5�_�   w   z           x           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �                 5�_�   x   {   y       z          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�     �               9        res=array.find_first with (item <15 & item >=13);5�_�   z   |           {      #    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�     �               A        res=array.find_first_index() with (item <15 & item >=13);5�_�   {   }           |      0    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�!     �               B        res=array.find_first_index(x) with (item <15 & item >=13);5�_�   |   ~           }      0    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�%     �               ?        res=array.find_first_index(x) with (x <15 & item >=13);5�_�   }              ~      -    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�+     �               =        res=array.find_first_index(x) with (x>5 & item >=13);5�_�   ~   �                 /    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�+     �               >        res=array.find_first_index(x) with (x >5 & item >=13);5�_�      �           �      =    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�.     �               ?        res=array.find_first_index(x) with (x > 5 & item >=13);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�=     �               (        $display("find_first : %p",res);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�J     �               9        res=array.find_first with (item <15 & item >=13);5�_�   �   �           �      *    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�^     �               8        res=array.find_last with (item <15 & item >=13);5�_�   �   �           �      6    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�g     �               8        res=array.find_last with (item <60 & item >=13);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�m     �               (        $display("find_first : %p",res);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�x     �               9        res=array.find_first with (item <15 & item >=13);5�_�   �   �           �      "    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�     �               @        res=array.find_last_index() with (item <15 & item >=13);5�_�   �   �           �      /    ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �               A        res=array.find_last_index(x) with (item <15 & item >=13);5�_�   �   �           �      0    ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �               >        res=array.find_last_index(x) with (x <15 & item >=13);5�_�   �   �           �      =    ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �               ?        res=array.find_last_index(x) with (x <100 & item >=13);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE��    �               (        $display("find_first : %p",res);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�.     �      	         %        $display("find(x) : %p",res);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�9     �   
            4        $display("find_index : res[%0d]=32",res[0]);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�C     �               (        $display("find_first : %p",res);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�K     �               .        $display("find_first item  : %p",res);5�_�   �   �           �      !    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�N     �               2        $display("find_first <=13item  : %p",res);5�_�   �   �           �      %    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�T     �               2        $display("find_first 13<=item  : %p",res);5�_�   �   �           �      #    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�\     �               .        $display("find_first_index : %p",res);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�m     �               '        $display("find_last : %p",res);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                 v        aE�x     �               ,        $display("find_last item : %p",res);5�_�   �   �           �      $    ����                                                                                                                                                                                                                                                                                                                                                 v        aE�    �               0        $display("find_last 20<=item : %p",res);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                            aF�'     �               
          5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                            aF�@     �                 $display("min :       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                            aF�E     �                 $display("The min :       5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                            aF�O     �               ,  $display("The minimum in array is :       5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                            aF�T     �               /  $display("The minimum in array %p is :       5�_�   �   �           �      *    ����                                                                                                                                                                                                                                                                                                                                                            aF�Y     �               0  $display("The minimum in array: %p is :       5�_�   �   �           �      3    ����                                                                                                                                                                                                                                                                                                                                                            aF�o     �               9  $display("The minimum in array: %p is : %p",array      5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                            aF�s     �               9  $display("The minimum in array: %p is : %p",array,res);5�_�   �   �           �      
    ����                                                                                                                                                                                                                                                                                                                                                            aF�v     �               A          $display("The minimum in array: %p is : %p",array,res);5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                            aF�y     �                5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                            aFą     �                       res = arrat.min();5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                                                            aFĊ     �                       vres = arrat.min();5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       aFē     �                        �             5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                v       aFĘ     �          "       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       aFĜ     �      #   "              �          "    5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                                                v       aFğ     �         %               res = arrat.min();5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                                                v       aFġ     �          %               res = arrat.min();5�_�   �   �           �      	    ����                                                                                                                                                                                                                                                                                                                                                v       aFı     �          %               res = arrat.min();5�_�   �   �           �   !        ����                                                                                                                                                                                                                                                                                                                                                v       aFĳ     �       #   %       5�_�   �   �           �   "        ����                                                                                                                                                                                                                                                                                                                                                v       aFĶ     �   !   &   &       �   "   #   &    5�_�   �   �           �   "        ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �   !   #   )       res = arrat.min();5�_�   �   �           �   "   	    ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �   !   #   )               res = arrat.min();5�_�   �   �           �   %        ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �   $   &   )       5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �   $   )   )              �   %   &   )    5�_�   �   �           �   %   	    ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �   $   &   ,               res = arrat.min();5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �         ,              res = arrat.min();5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �         ,      ?        $display("The minimum in array: %p is : %p",array,res);5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �         ,      -        $display("find_last_index : %p",res);5�_�   �   �           �      2    ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �         ,      ?        $display("The minimum in array: %p is : %p",array,res);5�_�   �   �           �      2    ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �         ,      ?        $display("The maximum in array: %p is : %p",array,res);5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       aF��     �          ,              res = arrat.min();5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       aF�	     �         ,              res = arrat.min();5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       aF�     �         ,              res = arrat.max();5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                v       aF�     �          ,              res = arrat.unique();5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                v       aF�     �   !   #   ,              res = arrat.min();5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                v       aF�     �      !   ,      ?        $display("The minimum in array: %p is : %p",array,res);5�_�   �   �           �       5    ����                                                                                                                                                                                                                                                                                                                                                v       aF�&     �      !   ,      G        $display("The unique memebers in array: %p is : %p",array,res);5�_�   �   �           �       3    ����                                                                                                                                                                                                                                                                                                                                                v       aF�)     �      !   ,      H        $display("The unique memebers in array: %p are : %p",array,res);5�_�   �   �           �      &    ����                                                                                                                                                                                                                                                                                                                                                v       aF�3     �         ,      /    int array[9]='{12,14,32,45,56,76,47,72,94};5�_�   �   �           �      (    ����                                                                                                                                                                                                                                                                                                                                                v       aF�4     �         ,      0    int array[9]='{12,14,32,45,56,76,4i7,72,94};5�_�   �   �           �      '    ����                                                                                                                                                                                                                                                                                                                                                v       aF�<     �         ,      /    int array[9]='{12,14,32,45,56,76,42,72,94};5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                v       aF�F     �   !   #   ,              res = array.min();5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                v       aF�J     �   !   #   ,              res = array.unique();5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                v       aF�N     �   !   #   ,              res = array.unique(x);5�_�   �   �           �   "   $    ����                                                                                                                                                                                                                                                                                                                                                v       aF�T     �   !   #   ,      &        res = array.unique(x) with ();5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                                v       aF�a     �   "   $   ,      ?        $display("The minimum in array: %p is : %p",array,res);5�_�   �   �           �   #   -    ����                                                                                                                                                                                                                                                                                                                                                v       aF�n     �   "   $   ,      F        $display("The unique members in array: %p is : %p",array,res);5�_�   �   �           �   #   .    ����                                                                                                                                                                                                                                                                                                                                                v       aF�q     �   "   $   ,      J        $display("The unique members in array <50: %p is : %p",array,res);5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                                                v       aFń     �   $   &   ,              res = arrat.min();5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                                                v       aFň     �   $   &   ,              res = array.min();5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                                v       aFŐ     �   %   '   ,      ?        $display("The minimum in array: %p is : %p",array,res);5�_�   �   �           �   '        ����                                                                                                                                                                                                                                                                                                                                                v       aFŧ     �   &   )   )      i       end�   &   (   *      i    �   &   (   +      i    �   &   (   ,      i    �   &   (   ,       5�_�   �   �           �   '        ����                                                                                                                                                                                                                                                                                                                                                v       aFū     �   %   '   )      O        $display("The index of unique members in array: %p is : %p",array,res);   i�   &   (   )      i5�_�   �   �           �   &   P    ����                                                                                                                                                                                                                                                                                                                                                v       aFŮ    �   %   )   (      P        $display("The index of unique members in array: %p is : %p",array,res);i5�_�   �   �           �   "   )    ����                                                                                                                                                                                                                                                                                                                                                v       aH�     �   !   #   *      *        res = array.unique(x) with (x<50);5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                v       aH�    �   !   #   *              res = array.unique(x);5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                                v       aH    �   !   #   *      !        res = array.unique(x<50);5�_�   �   �           �       !    ����                                                                                                                                                                                                                                                                                                                                                v       aH9     �      !   *      K        $display("The unique memebers in array: %p is/are : %p",array,res);5�_�   �   �           �   #   .    ����                                                                                                                                                                                                                                                                                                                                                v       aH@     �   "   $   *      U        $display("The unique members in array with value <50: %p is : %p",array,res);5�_�   �   �           �   #   D    ����                                                                                                                                                                                                                                                                                                                                                v       aHF     �   "   $   *      X        $display("The unique members in array %p with value <50: %p is : %p",array,res);5�_�   �   �           �   #   C    ����                                                                                                                                                                                                                                                                                                                                                v       aHK     �   "   $   *      T        $display("The unique members in array %p with value <50 is : %p",array,res);5�_�   �   �           �   #   D    ����                                                                                                                                                                                                                                                                                                                                                v       aHN   	 �   "   $   *      T        $display("The unique members in array %p with value <50 are: %p",array,res);5�_�   �   �           �   %       ����                                                                                                                                                                                                                                                                                                                                                v       aL     �   $   &   *      #        res = array.unique_index();5�_�   �   �           �   '        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL     �   &   )   *       5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL     �   '   ,   +       �   (   )   +    5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL     �   '   )   .       res = array.unique_index();5�_�   �   �           �   (   
    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL      �   '   )   .      %        i res = array.unique_index();5�_�   �   �           �   (        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL)     �   '   )   .      #        res = array.unique_index();5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL?     �   '   )   .              res = array.reverse();5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL@     �   '   )   .              res = array.reverse();i5�_�   �   �           �   )   6    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLJ     �   (   *   .      O        $display("The index of unique members in array: %p is : %p",array,res);5�_�   �   �           �   )       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL_   
 �   (   *   .      2        $display("reverse: %p is : %p",array,res);5�_�   �   �           �   +        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   *   /   .       �   +   ,   .    5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   .   3   1       �   /   0   1    5�_�   �   �           �   2        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   1   6   4       �   2   3   4    5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   *   ,   7       res = array.unique_index();5�_�   �   �           �   +        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   *   ,   7      #        res = array.unique_index();5�_�   �   �           �   -        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   ,   .   7       5�_�   �   �           �   -       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   ,   .   7      i5�_�   �   �           �   ,   I    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   +   -   7      O        $display("The index of unique members in array: %p is : %p",array,res);5�_�   �   �           �   ,   ?    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL     �   +   -   7      I        $display("The index of unique members in array: %p is : %p",res);5�_�   �   �           �   /       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL     �   .   0   7       res = array.unique_index();5�_�   �   �           �   /        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL     �   .   0   7      #        res = array.unique_index();5�_�   �   �           �   0   J    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL'     �   /   1   7      O        $display("The index of unique members in array: %p is : %p",array,res);5�_�   �   �           �   2        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL;     �   1   3   7       res = array.unique_index();5�_�   �   �           �   2   	    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL=     �   1   3   7      $         res = array.unique_index();5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLD     �   1   4   7      #        res = array.unique_index();5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLE     �   1   3   8              5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLH     �   1   3   8              for ()5�_�   �   �           �   2       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLS     �   2   4   9                     #        res = array.unique_index();�   1   4   8              for (int i=0;i<5;i++)5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLc     �   2   4   8      '            res = array.unique_index();5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLf     �   2   4   8      '            resi= array.unique_index();5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLh     �   2   4   8      '            resi= array.unique_index();5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLq     �   2   4   8      '            resi= array.unique_index();5�_�   �   �           �   3       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aLv     �   2   4   8      !            array.unique_index();5�_�   �   �           �   4   >    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   3   5   8      O        $display("The index of unique members in array: %p is : %p",array,res);5�_�   �   �           �   4   +    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   3   5   8      ;        $display("shuffle iteration:%0d = : %p",array,res);5�_�   �   �           �   4   7    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   3   5   8      9        $display("shuffle iteration:%0d = %p",array,res);5�_�   �   �           �   4   .    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   3   5   8      5        $display("shuffle iteration:%0d = %p",array);5�_�   �   �           �   4       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   3   5   8      7        $display("shuffle iteration:%0d = %p",i,array);5�_�   �   �           �   5        ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�    �   4   6   8       5�_�   �   �           �   (       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   '   )   8              res = array.reverse();5�_�   �   �           �   )   "    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�    �   (   *   8      $        $display("reverse: %p",res);5�_�   �   �           �   +       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   *   ,   8              res = array.sort();5�_�   �   �           �   ,       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   +   -   8      #        $display("sort =  %p",res);5�_�   �              �   ,   !    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   +   -   8      #        $display("sort =  %p",res);5�_�   �                /       ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL�     �   .   0   8              res = array.rsort();5�_�                    0   "    ����                                                                                                                                                                                                                                                                                                                           %          '           v       aL     �   /   1   8      $        $display("rsort =  %p",res);5�_�   x           z   y           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �              5�_�   q           s   r           ����                                                                                                                                                                                                                                                                                                                                                 v        aE��     �             �                          9        res=array.find_first with (item <15 & item >=13);   (        $display("find_first : %p",res);   
                  5�_�   &           (   '           ����                                                                                                                                                                                                                                                                                                                                                            aE��     �               m5��