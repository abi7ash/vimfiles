Vim�UnDo� �zF�Z"��J)����Awѽ��������    4   +        $display("xor   =%0h",array.xor());   2         j       j   j   j    aP�}   	 _�                             ����                                                                                                                                                                                                                                                                                                                                                             aO9&     �          8      
module tb;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             aO9'     �          9       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             aO9(     �          :       5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             aO9.     �          ;       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aO9Z     �         @          function new()5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aO9[     �         @          function new ()5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aO9^     �         @          function new (string name)5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                             aO9{     �   
      E              $display();5�_�      
           	      -    ����                                                                                                                                                                                                                                                                                                                                                             aO9�     �   
      E      /        $display(""name=%s rank=%0d pages=%0d);5�_�   	              
      ?    ����                                                                                                                                                                                                                                                                                                                                                             aO9�     �         I           �   
      E      ?        $display(""name=%s rank=%0d pages=%0d,name,rank,pages);5�_�   
                         ����                                                                                                                                                                                                                                                                                                                                                             aO9�     �         H      /    int array[9]='{12,14,32,45,56,76,45,72,94};5�_�                            ����                                                                                                                                                                                                                                                                                                                                       F           v       aO9�     �         H   5   /    int array[9]='{12,14,32,45,56,76,45,72,94};       int res[$];           initial begin   %        res=array.find(x) with (x>3);   '        $display("find(x>3) : %p",res);       /        res=array.find_index with (item == 32);   :        $display("find_index of 32 : res[%0d]=32",res[0]);       9        res=array.find_first with (item <15 & item >=13);   5        $display("find_first 13<=item<15  : %p",res);              3        res=array.find_first_index(x) with (x > 5);   8        $display("find_first_index for item>5: %p",res);   	            8        res=array.find_last with (item <60 & item >=20);   3        $display("find_last 20<=item<60 : %p",res);   	            3        res=array.find_last_index(x) with (x <100);   /        $display("find_last_index : %p\n",res);                  res = array.min();   A        $display("The minimum in array: %p is : %p\n",array,res);               res = array.max();   A        $display("The maximum in array: %p is : %p\n",array,res);               res = array.unique();   J        $display("The unique members in array: %p is/are : %p",array,res);       *        res = array.unique(x) with (x<50);   T        $display("The unique members in array %p with value <50 are: %p",array,res);       #        res = array.unique_index();   O        $display("The index of unique members in array: %p is : %p",array,res);               array.reverse();   &        $display("reverse: %p",array);               array.sort();   %        $display("sort =  %p",array);                   array.rsort();   &        $display("rsort =  %p",array);       #        for (int i=0;i<5;i++) begin               array.shuffle();   ;            $display("shuffle iteration:%0d = %p",i,array);           end           end5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aO9�     �                   5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                  v       aO9�     �                   initla begin5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aO9�     �                   5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v       aO9�     �                   5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v       aO9�     �               string n    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aO9�     �                   string n    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aO:     �               !    string name_arr[4] = '{};    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aO:     �               #    string name_arr[4] = '{""};    5�_�                       "    ����                                                                                                                                                                                                                                                                                                                                                  v       aO:	     �               (    string name_arr[4] = '{"alexa"};    5�_�                       $    ����                                                                                                                                                                                                                                                                                                                                                  v       aO:     �               +    string name_arr[4] = '{"alexa",""};    5�_�                       )    ����                                                                                                                                                                                                                                                                                                                                                  v       aO:     �               /    string name_arr[4] = '{"alexa","siri"};    5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                                  v       aO:     �               2    string name_arr[4] = '{"alexa","siri",""};    5�_�                       7    ����                                                                                                                                                                                                                                                                                                                                                  v       aO:     �               =    string name_arr[4] = '{"alexa","siri","google home"};    5�_�                       9    ����                                                                                                                                                                                                                                                                                                                                                  v       aO:     �               @    string name_arr[4] = '{"alexa","siri","google home",""};    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v       aO:      �                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aO:@     �               -----------Initial Values5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aO:A     �               ----------- Initial Values5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aO:T     �                       foreach()5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v       aO:_     �                       foreach(rt[i])5�_�      !                       ����                                                                                                                                                                                                                                                                                                                                                  v       aO:f     �               foreach(rt[i]) begin5�_�       "           !           ����                                                                                                                                                                                                                                                                                                                                                  v       aO:i     �                5�_�   !   #           "           ����                                                                                                                                                                                                                                                                                                                                                  v        aO:�     �      (           �              5�_�   "   $           #   &        ����                                                                                                                                                                                                                                                                                                                                                  v        aO:�     �   %   0   )       �   &   '   )    5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                  v        aO:�     �          2      )----------- Initial Values -----------");5�_�   $   &           %           ����                                                                                                                                                                                                                                                                                                                                                  v        aO:�     �      "   2              foreach(rt[i]) begin5�_�   %   '           &           ����                                                                                                                                                                                                                                                                                                                                                  v        aO:�     �      !   3              5�_�   &   (           '           ����                                                                                                                                                                                                                                                                                                                                                  v        aO:�     �      !   3              rt.sort()5�_�   '   )           (           ����                                                                                                                                                                                                                                                                                                                                                  v        aO:�     �      !   3              rt.sort(x)5�_�   (   +           )   !       ����                                                                                                                                                                                                                                                                                                                                                  v        aO:�     �       "   3              foreach(rt[i]) begin5�_�   )   ,   *       +   "       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;     �   !   "          &            rt[i] = new (name_arr[i]);5�_�   +   -           ,   "       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;     �   !   "                      rt[i].randomize();5�_�   ,   .           -   #       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;     �   "   #                  end5�_�   -   /           .   %       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;     �   $   &   0      )----------- Initial Values -----------");5�_�   .   0           /   &       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;4     �   %   (   0              foreach(rt[i]) begin5�_�   /   1           0   &       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;:     �   %   '   1              5�_�   0   2           1   (   &    ����                                                                                                                                                                                                                                                                                                                                                  v        aO;g     �   '   )   1      &            rt[i] = new (name_arr[i]);5�_�   1   3           2   (       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;j     �   '   (          &            rt[i] = new (name_arr[i]);5�_�   2   4           3   (       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;k     �   '   (                      rt[i].randomize();5�_�   3   5           4   )       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;o     �   (   *   /              end5�_�   4   6           5   )       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;v     �   (   *   /              5�_�   5   7           6   )       ����                                                                                                                                                                                                                                                                                                                                                  v        aO;x     �   (   )                  5�_�   6   8           7   )        ����                                                                                                                                                                                                                                                                                                                                                  v        aO;y     �   (   )           5�_�   7   9           8   )        ����                                                                                                                                                                                                                                                                                                                                                  v        aO;y     �   (   )           5�_�   8   ;           9   )        ����                                                                                                                                                                                                                                                                                                                                                  v        aO;z    �   (   )           5�_�   9   <   :       ;          ����                                                                                                                                                                                                                                                                                                                                                  v        aO;�     �   
      +      ?        $display(""name=%s rank=%0d pages=%0d,name,rank,pages);5�_�   ;   =           <      ,    ����                                                                                                                                                                                                                                                                                                                                                  v        aO;�     �   
      +      >        $display("name=%s rank=%0d pages=%0d,name,rank,pages);5�_�   <   ?           =      .    ����                                                                                                                                                                                                                                                                                                                                                  v        aO;�    �   
      +      @        $display("name=%s rank=%0d pages=%0d":,name,rank,pages);5�_�   =   @   >       ?          ����                                                                                                                                                                                                                                                                                                                                                  v        aO<     �         +              $display("   )----------- Initial Values -----------");�         +              $display("5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                  v        aO<!     �         *              $display("   '----------- Sort by name -----------");�         *              $display("5�_�   @   B           A   "       ����                                                                                                                                                                                                                                                                                                                                                  v        aO<$    �   !   #   )              $display("   .----------- Sort by rank, pages -----------");�   !   #   )              $display("5�_�   A   C           B   $       ����                                                                                                                                                                                                                                                                                                                                                  v        aP�2    �   #   %   (              foreach(rt[i]) begin5�_�   B   D           C           ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �         (       5�_�   C   E           D           ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �         )       5�_�   D   F           E   )        ����                                                                                                                                                                                                                                                                                                                                                   v        aP�     �   (   -   +       5�_�   E   G           F   +        ����                                                                                                                                                                                                                                                                                                                                                   v        aP�#     �   *   ,   .       5�_�   F   H           G   ,       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�.     �   +   -   .              $display()5�_�   G   I           H   ,       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�1     �   +   -   .              $display();5�_�   H   J           I   ,       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�>     �   +   -   .      !        $display("",array.sum());5�_�   I   L           J   -       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�[     �   ,   .   .          end5�_�   J   M   K       L   -       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�a     �   ,   /   .          end5�_�   L   N           M   -       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�c     �   -   0   /    �   -   .   /    5�_�   M   O           N   .       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�i     �   .   1   1    �   .   /   1    5�_�   N   P           O   /       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�m     �   /   2   3    �   /   0   3    5�_�   O   Q           P   0       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�n     �   0   3   5    �   0   1   5    5�_�   P   R           Q   .       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�}     �   -   /   7      +        $display("sum   =%0d",array.sum());5�_�   Q   S           R   .       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   -   /   7      0        $display("prroduct   =%0d",array.sum());5�_�   R   T           S   .   )    ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   -   /   7      -        $display("prroduct=%0d",array.sum());5�_�   S   U           T   /   '    ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   .   0   7      +        $display("sum   =%0d",array.sum());5�_�   T   V           U   /   &    ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   .   0   7      ,        $display("sum   =%0d",array.adnd());5�_�   U   W           V   0   '    ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   /   1   7      +        $display("sum   =%0d",array.sum());5�_�   V   X           W   1   '    ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   0   2   7      +        $display("sum   =%0d",array.sum());5�_�   W   Y           X   1       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   0   2   7      +        $display("sum   =%0d",array.xor());5�_�   X   Z           Y   0       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   /   1   7      *        $display("sum   =%0d",array.or());5�_�   Y   [           Z   /       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   .   0   7      +        $display("sum   =%0d",array.and());5�_�   Z   \           [   2       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   1   2              end5�_�   [   ]           \   2       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   1   2              end5�_�   \   ^           ]   2       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   1   2              end5�_�   ]   _           ^   2       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��    �   1   2              end5�_�   ^   `           _   +   !    ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   *   -   3      !        //Array reduction methods5�_�   _   a           `   ,       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   +   -   4              $display()5�_�   `   b           a   ,   $    ����                                                                                                                                                                                                                                                                                                                                                   v        aP��     �   +   -   4      $        $display(array  = %p",array)5�_�   a   c           b   ,       ����                                                                                                                                                                                                                                                                                                                                                   v        aP��    �   +   -   4      %        $display(array  = %p",array);5�_�   b   d           c   0       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�F     �   /   1   4      +        $display("and   =%0d",array.and());5�_�   c   e           d   0       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�O     �   /   1   4      *        $display("and   =%h",array.and());5�_�   d   f           e   1       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�Q     �   0   2   4      )        $display("or   =%0d",array.or());5�_�   e   g           f   2       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�T    �   1   3   4      +        $display("xor   =%0d",array.xor());5�_�   f   h           g   0        ����                                                                                                                                                                                                                                                                                                                                                   v        aP�j     �   /   1   4      +        $display("and   =%0h",array.and());5�_�   g   i           h   0       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�s     �   /   1   4      *       $display("and   =%0h",array.and());5�_�   h   j           i   1       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�y     �   0   2   4      )        $display("or   =%0h",array.or());5�_�   i               j   2       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�|   	 �   1   3   4      +        $display("xor   =%0h",array.xor());5�_�   J           L   K   -       ����                                                                                                                                                                                                                                                                                                                                                   v        aP�]     �   -   .   .    �   -   .   .      +        $display("sum   =%0d",array.sum());       end5�_�   =           ?   >          ����                                                                                                                                                                                                                                                                                                                                                  v        aO<     �         +              $display"5�_�   9           ;   :          ����                                                                                                                                                                                                                                                                                                                                                  v        aO;�     �   
           5�_�   )           +   *   !       ����                                                                                                                                                                                                                                                                                                                                                  v        aO:�     �       "        5��