Vim�UnDo� ?@�5*�<\�������U �ڐ�{��i   !   7                    6:"betray",8:"brazzen",21:"brink"};      5     �      �  �  �    aD��   	 _�                             ����                                                                                                                                                                                                                                                                                                                                       9   	       v   	    aD�~     �               9   
module tb;       (    //create a dynamic array of type int       int array[];       $    //dynamic array to hold a string       string fruits[];       5    //create a new array id and replicate it to array       int id[];           initial begin   /        //create dynamic array to hold 5 values           array = new[5];       /        //initialize the array with five values           foreach(array[i]) begin               array[i]=0;   ;            $display("clearing array[%0d]=%0d",i,array[i]);   H            array[i]=($random%100<0) ?(-1*($random%100)) : $random%100 ;   Y            $display("Adding a random value less than 100 to array[%0d]=%0d",i,array[i]);           end       %        //print the contents of array   %        $display("array = %p",array);   �        $display("\nLooks like tha value generated is not random...\nit seems to add the same value in each run..!!!\n:array = '{-99, 9, 57, 14, 29}\n ");          A        //create a dynamic array that can hold a string of values           fruits=new[3];              1        //initialize fruits with a set of strings   -        fruits = '{"apple","orange","mango"};   /        $display("\n \n fruits=%p\n\n",fruits);       %        //print the size of the array   8        $display("size of fruits is %0d",fruits.size());       *        //delete the contents of the array           fruits.delete();   X        $display("\n\nAfter doing fuits.delete(), fruits.size()=%0d\n\n",fruits.size());       '        //replicate id to contain array           id = array;                      //show contents of id   k        $display("\narray contents have been replicated to id.\nso id=%p and size of id=%0d",id,id.size());       +        //add another another element to id   "        id = new[id.size()+1](id);           id[id.size()-1]=6;       *        //compare contents of id and array   Z        $display("\nnow added a new element '6' to id alone.\nid=%p \narray=%p",id,array);           end       	endmodule5�_�                            ����                                                                                                                                                                                                                                                                                                                                          	       v   	    aDڄ     �                   5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                       
   	       v   	    aDډ     �         
                       1                                   "orange" : 10,�         	      *              fruits_l0 = '{ "apple"  : 4,5�_�                       *    ����                                                                                                                                                                                                                                                                                                                                       
   	       v   	    aDڑ     �         	      *              fruits_l0 = '{ "apple"  : 4,   >                                                "orange" : 10,�         	      *              fruits_l0 = '{ "apple"  : 4,5�_�                       8    ����                                                                                                                                                                                                                                                                                                                                       	   	       v   	    aDژ     �               8              fruits_l0 = '{ "apple"  : 4,"orange" : 10,   E                                                        "plum"   : 9,�               8              fruits_l0 = '{ "apple"  : 4,"orange" : 10,5�_�                       E    ����                                                                                                                                                                                                                                                                                                                                          	       v   	    aDڝ     �               E              fruits_l0 = '{ "apple"  : 4,"orange" : 10,"plum"   : 9,   \                                                                             "guava"  : 1 };�               E              fruits_l0 = '{ "apple"  : 4,"orange" : 10,"plum"   : 9,5�_�      
                 T    ����                                                                                                                                                                                                                                                                                                                                          	       v   	    aDڧ     �      $         T              fruits_l0 = '{ "apple"  : 4,"orange" : 10,"plum"   : 9,"guava"  : 1 };5�_�                
          ����                                                                                                                                                                                                                                                                                                                                       %   	       v   	    aD��     �         $      S                   // size() : Print the number of items in the given dynamic array5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD��     �      	   %      O                         $display ("fruits_l0.size() = %0d", fruits_l0.size());5�_�                           ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD��     �   
      %      b                               // num() : Another function to print number of items in given array5�_�                       %    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD��     �         %      Y                                     $display ("fruits_l0.num() = %0d", fruits_l0.num());5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      o                                           // exists() : Check if a particular key exists in this dynamic array5�_�                       1    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      Q                                                 if (fruits_l0.exists ("orange"))5�_�                       =    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      r                                                             $display ("Found %0d orange !", fruits_l0["orange"]);5�_�                       C    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      f                                                                   if (!fruits_l0.exists ("apricots"))5�_�                       O    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      �                                                                               $display ("Sorry, season for apricots is over ...");5�_�                       U    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�&     �         %      �                                                                                     // Note: String indices are taken in alphabetical order5�_�                           ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      �                                                                                           // first() : Get the first element in the array5�_�                           ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      �                                                                                           // first() : Get the first element in the array5�_�                       W    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      �                                                                                       // first() : Get the first element in the array5�_�                       S    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      �                                                                                   // first() : Get the first element in the array5�_�                       O    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      ~                                                                               // first() : Get the first element in the array5�_�                       K    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      z                                                                           // first() : Get the first element in the array5�_�                       G    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      v                                                                       // first() : Get the first element in the array5�_�                       C    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      r                                                                   // first() : Get the first element in the array5�_�                       ?    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      n                                                               // first() : Get the first element in the array5�_�                       ;    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      j                                                           // first() : Get the first element in the array5�_�                       7    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      f                                                       // first() : Get the first element in the array5�_�                        3    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      b                                                   // first() : Get the first element in the array5�_�      !                  /    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      ^                                               // first() : Get the first element in the array5�_�       "           !      +    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      Z                                           // first() : Get the first element in the array5�_�   !   #           "      '    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      V                                       // first() : Get the first element in the array5�_�   "   $           #      #    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      R                                   // first() : Get the first element in the array5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      N                               // first() : Get the first element in the array5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      J                           // first() : Get the first element in the array5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      F                       // first() : Get the first element in the array5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�     �         %      B                   // first() : Get the first element in the array5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�#     �         %      f                                                                                                 begin5�_�   (   *           )      ]    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�$     �         %      b                                                                                             begin5�_�   )   +           *      Y    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�$     �         %      ^                                                                                         begin5�_�   *   ,           +      U    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�$     �         %      Z                                                                                     begin5�_�   +   -           ,      Q    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�$     �         %      V                                                                                 begin5�_�   ,   .           -      M    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�$     �         %      R                                                                             begin5�_�   -   /           .      I    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�$     �         %      N                                                                         begin5�_�   .   0           /      E    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�$     �         %      J                                                                     begin5�_�   /   1           0      A    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�$     �         %      F                                                                 begin5�_�   0   2           1      =    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�$     �         %      B                                                             begin5�_�   1   3           2      9    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�%     �         %      >                                                         begin5�_�   2   4           3      5    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�%     �         %      :                                                     begin5�_�   3   5           4      1    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�%     �         %      6                                                 begin5�_�   4   6           5      -    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�%     �         %      2                                             begin5�_�   5   7           6      )    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�&     �         %      .                                         begin5�_�   6   8           7      %    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�&     �         %      *                                     begin5�_�   7   9           8      !    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�'     �         %      &                                 begin5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�'     �         %      "                             begin5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�(     �         %                               begin5�_�   :   <           ;          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�(     �         %                           begin5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�,     �         %                       begin5�_�   <   >           =          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�D     �         %      r                                                                                                         string f;5�_�   =   ?           >      e    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�D     �         %      n                                                                                                     string f;5�_�   >   @           ?      a    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�D     �         %      j                                                                                                 string f;5�_�   ?   A           @      ]    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�D     �         %      f                                                                                             string f;5�_�   @   B           A      Y    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�D     �         %      b                                                                                         string f;5�_�   A   C           B      U    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�E     �         %      ^                                                                                     string f;5�_�   B   D           C      Q    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�E     �         %      Z                                                                                 string f;5�_�   C   E           D      M    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�E     �         %      V                                                                             string f;5�_�   D   F           E      I    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�E     �         %      R                                                                         string f;5�_�   E   G           F      E    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�E     �         %      N                                                                     string f;5�_�   F   H           G      A    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�E     �         %      J                                                                 string f;5�_�   G   I           H      =    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�E     �         %      F                                                             string f;5�_�   H   J           I      9    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�F     �         %      B                                                         string f;5�_�   I   K           J      5    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�F     �         %      >                                                     string f;5�_�   J   L           K      1    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�F     �         %      :                                                 string f;5�_�   K   M           L      -    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�F     �         %      6                                             string f;5�_�   L   N           M      )    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�F     �         %      2                                         string f;5�_�   M   O           N      %    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�G     �         %      .                                     string f;5�_�   N   P           O      !    ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�G     �         %      *                                 string f;5�_�   O   Q           P          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�H     �         %      &                             string f;5�_�   P   R           Q          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�H     �         %      "                         string f;5�_�   Q   S           R          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�I     �         %                           string f;5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�J     �         %                       string f;5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD�n     �         %                   begin5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                                       '   	       v   	    aD�q     �         &                   5�_�   U   W           V           ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܃     �          *      �                                                                                                                 // This function returns true if it succeeded and first key is stored5�_�   V   X           W           ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܈     �          *      �                                                                                                                 // This function returns true if it succeeded and first key is stored5�_�   W   Y           X      m    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܈     �          *      �                                                                                                             // This function returns true if it succeeded and first key is stored5�_�   X   Z           Y      i    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܈     �          *      �                                                                                                         // This function returns true if it succeeded and first key is stored5�_�   Y   [           Z      e    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܈     �          *      �                                                                                                     // This function returns true if it succeeded and first key is stored5�_�   Z   \           [      a    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܈     �          *      �                                                                                                 // This function returns true if it succeeded and first key is stored5�_�   [   ]           \      ]    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܈     �          *      �                                                                                             // This function returns true if it succeeded and first key is stored5�_�   \   ^           ]      Y    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܉     �          *      �                                                                                         // This function returns true if it succeeded and first key is stored5�_�   ]   _           ^      U    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܉     �          *      �                                                                                     // This function returns true if it succeeded and first key is stored5�_�   ^   `           _      Q    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܉     �          *      �                                                                                 // This function returns true if it succeeded and first key is stored5�_�   _   a           `      M    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܉     �          *      �                                                                             // This function returns true if it succeeded and first key is stored5�_�   `   b           a      I    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܊     �          *      �                                                                         // This function returns true if it succeeded and first key is stored5�_�   a   c           b      E    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܊     �          *      �                                                                     // This function returns true if it succeeded and first key is stored5�_�   b   d           c      A    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܊     �          *      �                                                                 // This function returns true if it succeeded and first key is stored5�_�   c   e           d      =    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܊     �          *      �                                                             // This function returns true if it succeeded and first key is stored5�_�   d   f           e      9    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܊     �          *      ~                                                         // This function returns true if it succeeded and first key is stored5�_�   e   g           f      5    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܊     �          *      z                                                     // This function returns true if it succeeded and first key is stored5�_�   f   h           g      1    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܊     �          *      v                                                 // This function returns true if it succeeded and first key is stored5�_�   g   i           h      -    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܋     �          *      r                                             // This function returns true if it succeeded and first key is stored5�_�   h   j           i      )    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܋     �          *      n                                         // This function returns true if it succeeded and first key is stored5�_�   i   k           j      %    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܌     �          *      j                                     // This function returns true if it succeeded and first key is stored5�_�   j   l           k      !    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܌     �          *      f                                 // This function returns true if it succeeded and first key is stored5�_�   k   m           l          ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܌     �          *      b                             // This function returns true if it succeeded and first key is stored5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܍     �          *      ^                         // This function returns true if it succeeded and first key is stored5�_�   m   o           n          ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܍     �          *      Z                     // This function returns true if it succeeded and first key is stored5�_�   n   p           o          ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܎     �          *      V                 // This function returns true if it succeeded and first key is stored5�_�   o   q           p          ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aD܏     �          *      R             // This function returns true if it succeeded and first key is stored5�_�   p   r           q      	    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܒ     �         *                   string f;5�_�   q   s           r      	    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܔ     �         *                   begin5�_�   r   t           s       	    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܘ     �      !   *      �                                                                                                                         // in the provided string "f"5�_�   s   u           t       u    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܘ     �      !   *      �                                                                                                                     // in the provided string "f"5�_�   t   v           u       q    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܘ     �      !   *      �                                                                                                                 // in the provided string "f"5�_�   u   w           v       m    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܘ     �      !   *      �                                                                                                             // in the provided string "f"5�_�   v   x           w       i    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      �                                                                                                         // in the provided string "f"5�_�   w   y           x       e    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      �                                                                                                     // in the provided string "f"5�_�   x   z           y       a    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      ~                                                                                                 // in the provided string "f"5�_�   y   {           z       ]    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      z                                                                                             // in the provided string "f"5�_�   z   |           {       Y    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      v                                                                                         // in the provided string "f"5�_�   {   }           |       U    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      r                                                                                     // in the provided string "f"5�_�   |   ~           }       Q    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      n                                                                                 // in the provided string "f"5�_�   }              ~       M    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      j                                                                             // in the provided string "f"5�_�   ~   �                  I    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      f                                                                         // in the provided string "f"5�_�      �           �       E    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      b                                                                     // in the provided string "f"5�_�   �   �           �       A    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      ^                                                                 // in the provided string "f"5�_�   �   �           �       =    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      Z                                                             // in the provided string "f"5�_�   �   �           �       9    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܙ     �      !   *      V                                                         // in the provided string "f"5�_�   �   �           �       5    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܚ     �      !   *      R                                                     // in the provided string "f"5�_�   �   �           �       1    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܚ     �      !   *      N                                                 // in the provided string "f"5�_�   �   �           �       -    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܚ     �      !   *      J                                             // in the provided string "f"5�_�   �   �           �       )    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܚ     �      !   *      F                                         // in the provided string "f"5�_�   �   �           �       %    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܚ     �      !   *      B                                     // in the provided string "f"5�_�   �   �           �       !    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܛ     �      !   *      >                                 // in the provided string "f"5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܛ     �      !   *      :                             // in the provided string "f"5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܛ     �      !   *      6                         // in the provided string "f"5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܛ     �      !   *      2                     // in the provided string "f"5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܜ     �      !   *      .                 // in the provided string "f"5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܜ     �      !   *      *             // in the provided string "f"5�_�   �   �           �   !   	    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      �                                                                                                                                 if (fruits_l0.first (f))5�_�   �   �           �   !   }    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      �                                                                                                                             if (fruits_l0.first (f))5�_�   �   �           �   !   y    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      �                                                                                                                         if (fruits_l0.first (f))5�_�   �   �           �   !   u    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      �                                                                                                                     if (fruits_l0.first (f))5�_�   �   �           �   !   q    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      �                                                                                                                 if (fruits_l0.first (f))5�_�   �   �           �   !   m    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      �                                                                                                             if (fruits_l0.first (f))5�_�   �   �           �   !   i    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      �                                                                                                         if (fruits_l0.first (f))5�_�   �   �           �   !   e    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      }                                                                                                     if (fruits_l0.first (f))5�_�   �   �           �   !   a    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      y                                                                                                 if (fruits_l0.first (f))5�_�   �   �           �   !   ]    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      u                                                                                             if (fruits_l0.first (f))5�_�   �   �           �   !   Y    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      q                                                                                         if (fruits_l0.first (f))5�_�   �   �           �   !   U    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      m                                                                                     if (fruits_l0.first (f))5�_�   �   �           �   !   Q    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܟ     �       "   *      i                                                                                 if (fruits_l0.first (f))5�_�   �   �           �   !   M    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      e                                                                             if (fruits_l0.first (f))5�_�   �   �           �   !   I    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      a                                                                         if (fruits_l0.first (f))5�_�   �   �           �   !   E    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      ]                                                                     if (fruits_l0.first (f))5�_�   �   �           �   !   A    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      Y                                                                 if (fruits_l0.first (f))5�_�   �   �           �   !   =    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      U                                                             if (fruits_l0.first (f))5�_�   �   �           �   !   9    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      Q                                                         if (fruits_l0.first (f))5�_�   �   �           �   !   5    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      M                                                     if (fruits_l0.first (f))5�_�   �   �           �   !   1    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      I                                                 if (fruits_l0.first (f))5�_�   �   �           �   !   -    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      E                                             if (fruits_l0.first (f))5�_�   �   �           �   !   )    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      A                                         if (fruits_l0.first (f))5�_�   �   �           �   !   %    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      =                                     if (fruits_l0.first (f))5�_�   �   �           �   !   !    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܠ     �       "   *      9                                 if (fruits_l0.first (f))5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܡ     �       "   *      5                             if (fruits_l0.first (f))5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܡ     �       "   *      1                         if (fruits_l0.first (f))5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܢ     �       "   *      -                     if (fruits_l0.first (f))5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܢ     �       "   *      )                 if (fruits_l0.first (f))5�_�   �   �           �   !       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܤ     �       "   *      %             if (fruits_l0.first (f))5�_�   �   �           �   "   �    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܧ     �   !   #   *      �                                                                                                                                               $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   �    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܧ     �   !   #   *      �                                                                                                                                           $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   �    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܧ     �   !   #   *      �                                                                                                                                       $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   �    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܧ     �   !   #   *      �                                                                                                                                   $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                                                               $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   {    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                                                           $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   w    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                                                       $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   s    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                                                   $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   o    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                                               $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   k    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                                           $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   g    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                                       $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   c    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                                   $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   _    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                               $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   [    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                           $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   W    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                       $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   S    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                                   $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   O    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                               $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   K    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                           $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   G    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      �                                                                       $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   C    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      |                                                                   $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   ?    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܨ     �   !   #   *      x                                                               $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   ;    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܩ     �   !   #   *      t                                                           $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   7    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܩ     �   !   #   *      p                                                       $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   3    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܩ     �   !   #   *      l                                                   $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   /    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܩ     �   !   #   *      h                                               $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   +    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܩ     �   !   #   *      d                                           $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   '    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܩ     �   !   #   *      `                                       $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "   #    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܩ     �   !   #   *      \                                   $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܩ     �   !   #   *      X                               $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܪ     �   !   #   *      T                           $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܫ     �   !   #   *      P                       $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܬ     �   !   #   *      L                   $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);5�_�   �   �           �   "       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܮ     �   !   $   *      H               $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);   �                                                                                                                                                     end5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܱ     �   "   $   *      �                                                                                                                                                 end5�_�   �   �           �   #   �    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܱ     �   "   $   *      �                                                                                                                                             end5�_�   �   �           �   #   �    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܱ     �   "   $   *      �                                                                                                                                         end5�_�   �   �           �   #   �    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܱ     �   "   $   *      �                                                                                                                                     end5�_�   �   �           �   #   �    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܱ     �   "   $   *      �                                                                                                                                 end5�_�   �   �           �   #   }    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܱ     �   "   $   *      �                                                                                                                             end5�_�   �   �           �   #   y    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܱ     �   "   $   *      |                                                                                                                         end5�_�   �   �           �   #   u    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܱ     �   "   $   *      x                                                                                                                     end5�_�   �   �           �   #   q    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܱ     �   "   $   *      t                                                                                                                 end5�_�   �   �           �   #   m    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      p                                                                                                             end5�_�   �   �           �   #   i    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      l                                                                                                         end5�_�   �   �           �   #   e    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      h                                                                                                     end5�_�   �   �           �   #   a    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      d                                                                                                 end5�_�   �   �           �   #   ]    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      `                                                                                             end5�_�   �   �           �   #   Y    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      \                                                                                         end5�_�   �   �           �   #   U    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      X                                                                                     end5�_�   �   �           �   #   Q    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      T                                                                                 end5�_�   �   �           �   #   M    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      P                                                                             end5�_�   �   �           �   #   I    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      L                                                                         end5�_�   �   �           �   #   E    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      H                                                                     end5�_�   �   �           �   #   A    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      D                                                                 end5�_�   �   �           �   #   =    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      @                                                             end5�_�   �   �           �   #   9    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      <                                                         end5�_�   �   �           �   #   5    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      8                                                     end5�_�   �   �           �   #   1    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܲ     �   "   $   *      4                                                 end5�_�   �   �           �   #   -    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܳ     �   "   $   *      0                                             end5�_�   �   �           �   #   )    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܳ     �   "   $   *      ,                                         end5�_�   �   �           �   #   %    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܳ     �   "   $   *      (                                     end5�_�   �   �           �   #   !    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܳ     �   "   $   *      $                                 end5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܳ     �   "   $   *                                    end5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܴ     �   "   $   *                               end5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܴ     �   "   $   *                           end5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܵ     �   "   $   *                       end5�_�   �   �           �   #       ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܶ     �   "   $   *                   end5�_�   �   �           �   #   	    ����                                                                                                                                                                                                                                                                                                                                       +   	       v   	    aDܸ     �   "   %   *               end5�_�   �   �   �       �   &   	    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                                                           // last() : Get the last element in the array5�_�   �   �           �   &   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                                                       // last() : Get the last element in the array5�_�   �   �           �   &   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                                                   // last() : Get the last element in the array5�_�   �   �           �   &   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                                               // last() : Get the last element in the array5�_�   �   �           �   &   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                                           // last() : Get the last element in the array5�_�   �   �           �   &   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                                       // last() : Get the last element in the array5�_�   �   �           �   &   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                                   // last() : Get the last element in the array5�_�   �   �           �   &       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                               // last() : Get the last element in the array5�_�   �   �           �   &   {    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                           // last() : Get the last element in the array5�_�   �   �           �   &   w    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                       // last() : Get the last element in the array5�_�   �   �           �   &   s    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                                   // last() : Get the last element in the array5�_�   �   �           �   &   o    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                               // last() : Get the last element in the array5�_�   �   �           �   &   k    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                           // last() : Get the last element in the array5�_�   �              �   &   g    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                       // last() : Get the last element in the array5�_�   �                &   c    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                                   // last() : Get the last element in the array5�_�                  &   _    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                               // last() : Get the last element in the array5�_�                 &   [    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                           // last() : Get the last element in the array5�_�                 &   W    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                       // last() : Get the last element in the array5�_�                 &   S    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      �                                                                                   // last() : Get the last element in the array5�_�                 &   O    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      |                                                                               // last() : Get the last element in the array5�_�                 &   K    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      x                                                                           // last() : Get the last element in the array5�_�                 &   G    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      t                                                                       // last() : Get the last element in the array5�_�    	             &   C    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      p                                                                   // last() : Get the last element in the array5�_�    
          	   &   ?    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      l                                                               // last() : Get the last element in the array5�_�  	            
   &   ;    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      h                                                           // last() : Get the last element in the array5�_�  
               &   7    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      d                                                       // last() : Get the last element in the array5�_�                 &   3    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      `                                                   // last() : Get the last element in the array5�_�                 &   /    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      \                                               // last() : Get the last element in the array5�_�                 &   +    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      X                                           // last() : Get the last element in the array5�_�                 &   '    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      T                                       // last() : Get the last element in the array5�_�                 &   #    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      P                                   // last() : Get the last element in the array5�_�                 &       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      L                               // last() : Get the last element in the array5�_�                 &       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      H                           // last() : Get the last element in the array5�_�                 &       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      D                       // last() : Get the last element in the array5�_�                 &       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      @                   // last() : Get the last element in the array5�_�                 &       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      <               // last() : Get the last element in the array5�_�                 &       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   %   '   +      8           // last() : Get the last element in the array5�_�                 '       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                                                                 begin5�_�                 '   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                                                             begin5�_�                 '   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                                                         begin5�_�                 '   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                                                     begin5�_�                 '   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                                                 begin5�_�                 '   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                                             begin5�_�                 '   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                                         begin5�_�                 '   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                                     begin5�_�                  '   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                                 begin5�_�    !              '   }    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      �                                                                                                                             begin5�_�     "          !   '   y    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      ~                                                                                                                         begin5�_�  !  #          "   '   u    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      z                                                                                                                     begin5�_�  "  $          #   '   q    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      v                                                                                                                 begin5�_�  #  %          $   '   m    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      r                                                                                                             begin5�_�  $  &          %   '   i    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      n                                                                                                         begin5�_�  %  '          &   '   e    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      j                                                                                                     begin5�_�  &  (          '   '   a    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      f                                                                                                 begin5�_�  '  )          (   '   ]    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      b                                                                                             begin5�_�  (  *          )   '   Y    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      ^                                                                                         begin5�_�  )  +          *   '   U    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      Z                                                                                     begin5�_�  *  ,          +   '   Q    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      V                                                                                 begin5�_�  +  -          ,   '   M    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      R                                                                             begin5�_�  ,  .          -   '   I    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      N                                                                         begin5�_�  -  /          .   '   E    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      J                                                                     begin5�_�  .  0          /   '   A    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      F                                                                 begin5�_�  /  1          0   '   =    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      B                                                             begin5�_�  0  2          1   '   9    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      >                                                         begin5�_�  1  3          2   '   5    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      :                                                     begin5�_�  2  4          3   '   1    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      6                                                 begin5�_�  3  5          4   '   -    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      2                                             begin5�_�  4  6          5   '   )    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      .                                         begin5�_�  5  7          6   '   %    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      *                                     begin5�_�  6  8          7   '   !    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      &                                 begin5�_�  7  9          8   '       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      "                             begin5�_�  8  :          9   '       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +                               begin5�_�  9  ;          :   '       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +                           begin5�_�  :  <          ;   '       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +                       begin5�_�  ;  =          <   '       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +                   begin5�_�  <  >          =   '   	    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +               begin5�_�  =  @          >   '       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   (   +      
     begin5�_�  >  A  ?      @   (       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                                                         string f;5�_�  @  B          A   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                                                     string f;5�_�  A  C          B   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                                                 string f;5�_�  B  D          C   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                                             string f;5�_�  C  E          D   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                                         string f;5�_�  D  F          E   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                                     string f;5�_�  E  G          F   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                                 string f;5�_�  F  H          G   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                             string f;5�_�  G  I          H   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                         string f;5�_�  H  J          I   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                     string f;5�_�  I  K          J   (   �    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                                 string f;5�_�  J  L          K   (   }    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                             string f;5�_�  K  M          L   (   y    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �                                                                                                                         string f;5�_�  L  N          M   (   u    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      ~                                                                                                                     string f;5�_�  M  O          N   (   q    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      z                                                                                                                 string f;5�_�  N  P          O   (   m    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      v                                                                                                             string f;5�_�  O  Q          P   (   i    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      r                                                                                                         string f;5�_�  P  R          Q   (   e    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      n                                                                                                     string f;5�_�  Q  S          R   (   a    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      j                                                                                                 string f;5�_�  R  T          S   (   ]    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      f                                                                                             string f;5�_�  S  U          T   (   Y    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      b                                                                                         string f;5�_�  T  V          U   (   U    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      ^                                                                                     string f;5�_�  U  W          V   (   Q    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      Z                                                                                 string f;5�_�  V  X          W   (   M    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      V                                                                             string f;5�_�  W  Y          X   (   I    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      R                                                                         string f;5�_�  X  Z          Y   (   E    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      N                                                                     string f;5�_�  Y  [          Z   (   A    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      J                                                                 string f;5�_�  Z  \          [   (   =    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      F                                                             string f;5�_�  [  ]          \   (   9    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      B                                                         string f;5�_�  \  ^          ]   (   5    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      >                                                     string f;5�_�  ]  _          ^   (   1    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      :                                                 string f;5�_�  ^  `          _   (   -    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      6                                             string f;5�_�  _  a          `   (   )    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      2                                         string f;5�_�  `  b          a   (   %    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      .                                     string f;5�_�  a  c          b   (   !    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      *                                 string f;5�_�  b  d          c   (       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      &                             string f;5�_�  c  e          d   (       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      "                         string f;5�_�  d  f          e   (       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +                           string f;5�_�  e  g          f   (       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +                       string f;5�_�  f  h          g   (       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +                   string f;5�_�  g  i          h   '   	    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   &   )   +              begin            string f;5�_�  h  j          i           ����                                                                                                                                                                                                                                                                                                                                       +           v        aD��     �              *        int      fruits_l0 [string];               initial begin   T              fruits_l0 = '{ "apple"  : 4,"orange" : 10,"plum"   : 9,"guava"  : 1 };                         P                // size() : Print the number of items in the given dynamic array   F                $display ("fruits_l0.size() = %0d", fruits_l0.size());           S                // num() : Another function to print number of items in given array   D                $display ("fruits_l0.num() = %0d", fruits_l0.num());           T                // exists() : Check if a particular key exists in this dynamic array   0                if (fruits_l0.exists ("orange"))   I                    $display ("Found %0d orange !", fruits_l0["orange"]);       3                if (!fruits_l0.exists ("apricots"))   H                    $display ("Sorry, season for apricots is over ...");       G                // Note: String indices are taken in alphabetical order   >               // first() : Get the first element in the array           end       	endmodule                    begin            string f;   N         // This function returns true if it succeeded and first key is stored   &         // in the provided string "f"   !         if (fruits_l0.first (f))   D           $display ("fruits_l0.first [%s] = %0d", f, fruits_l0[f]);   	                     end       4       // last() : Get the last element in the array   	    begin        string f;   �                                                                                                                                                                                 if (fruits_l0.last (f))   �                                                                                                                                                                                     -- p    5�_�  i  k          j           ����                                                                                                                                                                                                                                                                                                                                                  v        aD��     �                  5�_�  j  l          k          ����                                                                                                                                                                                                                                                                                                                                                  v        aD߆     �                             $display()5�_�  k  m          l           ����                                                                                                                                                                                                                                                                                                                                                  v        aDߒ     �                 "            $display(array1=%p,())5�_�  l  n          m      3    ����                                                                                                                                                                                                                                                                                                                                                  v        aD߫     �                 3            $display(array1=%p,(array1[i]=$random))5�_�  m  o          n           ����                                                                                                                                                                                                                                                                                                                                                  v        aD߽     �               4            $display(array1=%p,(array1[i]=$random));5�_�  n  p          o          ����                                                                                                                                                                                                                                                                                                                                                  v        aD��     �                            array1[i]=$random));5�_�  o  q          p          ����                                                                                                                                                                                                                                                                                                                                                  v        aD��     �                           array1[i]=$random;5�_�  p  r          q           ����                                                                                                                                                                                                                                                                                                                                                 v       aD��     �                �             5�_�  q  s          r           ����                                                                                                                                                                                                                                                                                                                                                 v       aD��     �                foreach(array1[i])5�_�  r  t          s          ����                                                                                                                                                                                                                                                                                                                                                 v       aD��     �                    foreach(array1[i])5�_�  s  u          t          ����                                                                                                                                                                                                                                                                                                                                                 v       aD��     �                        foreach(array1[i])5�_�  t  v          u      	    ����                                                                                                                                                                                                                                                                                                                                                 v       aD��     �               	        i5�_�  u  w          v          ����                                                                                                                                                                                                                                                                                                                                                 v       aD�      �                       foreach(array1[i])5�_�  v  x          w          ����                                                                                                                                                                                                                                                                                                                                                 v       aD�     �                           array1[i]=$random;5�_�  w  y          x          ����                                                                                                                                                                                                                                                                                                                                                 v       aD�     �                        $display("array1[i]=%p);5�_�  x  z          y           ����                                                                                                                                                                                                                                                                                                                                                 v       aD�     �                        $display("array2[i]=%p);5�_�  y  {          z           ����                                                                                                                                                                                                                                                                                                                                                 v       aD�      �                �             5�_�  z  |          {           ����                                                                                                                                                                                                                                                                                                                                                 v       aD�"     �                 foreach(array1[i])5�_�  {  }          |      	    ����                                                                                                                                                                                                                                                                                                                                                 v       aD�%     �                         foreach(array1[i])5�_�  |  ~          }          ����                                                                                                                                                                                                                                                                                                                                                 v       aD�+     �                        foreach(array1[i])5�_�  }            ~          ����                                                                                                                                                                                                                                                                                                                                                 v       aD�/     �                            array1[i]=$random;5�_�  ~  �                    ����                                                                                                                                                                                                                                                                                                                                                 v       aD�4     �                         $display("array1[i]=%p);5�_�    �          �           ����                                                                                                                                                                                                                                                                                                                                                 v       aD�9     �                         $display("array3[i]=%p);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                 v       aD�B    �         "          endmodule5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                                 v       aD�3     �   
      "       5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                 v       aD�6     �   
      "      i5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                v       aD�Q     �         "              foreach(array1[i])               array1[i]=$random;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�Z     �         !                 array1[i]=$random;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�^     �         !              array1[i]=$random;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�y     �         !              array1='{;5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD��     �         "      "                 7:22,9:33,24:54};5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD��     �         "               $display("array1[i]=%p);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD��     �         "              $display("array1=%p);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "              foreach(array2[i])5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "          5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "         5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "        5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�      �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�!     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�"     �         "       5�_�  �  �          �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�'     �         "                      array2[i]=$random;�         "       5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�4     �         !              array2[i]=$random;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�N     �         !              array2[i]='{2:"";5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�X     �         !              array2[i]='{2:"beauty";5�_�  �  �  �      �          ����                                                                                                                                                                                                                                                                                                                                         
       v       aD��     �         "               $display("array2[i]=%p);5�_�  �  �  �      �           ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �                        foreach(array3[i])5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !                  array3[i]=$random;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !      2        array2[i]='{2:"beauty",4:"baker",5:"bitch"5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !              array3[i]=$random;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !              array3=$random;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD��     �         !      (        array3='{a:"tamil",b:"korean",d;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD��     �         !      )        array3='{"a:"tamil",b:"korean",d;5�_�  �  �          �   
       ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �   	      !              array3=new[6];5�_�  �  �          �      *    ����                                                                                                                                                                                                                                                                                                                                                V       aD�      �         !      *        array3='{"a":"tamil",b:"korean",d;5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�(     �         !               $display("array3[i]=%p);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�,     �         !              $display("array3=%p);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�;    �         !              $display("array1=%p");5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�4     �         !              array1='{1:32,2:23,4:435�_�  �  �          �      /    ����                                                                                                                                                                                                                                                                                                                                                V       aD�=    �         !      /        array2='{2:"beauty",4:"baker",5:"bitch"5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�s     �         !      )        array3='{"a":"tamil",b:"korean");5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�w    �         !      *        array3='{"a":"tamil","b:"korean");5�_�  �  �          �      *    ����                                                                                                                                                                                                                                                                                                                                                V       aD�    �         !      +        array3='{"a":"tamil","b":"korean");5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD��    �         !          string arrat3[string];5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD��     �      	   !              array1=new[5];5�_�  �  �          �   	       ����                                                                                                                                                                                                                                                                                                                                                V       aD��     �      
   !              array2=new[4];5�_�  �  �          �   
       ����                                                                                                                                                                                                                                                                                                                                                V       aD��    �   	      !              array3=new[2];5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !      (        $display("array2[i]=%p",array2);5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !      0        array2='{2:"beauty",4:"baker",5:"bitch",5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !      .        array2='{"beauty",4:"baker",5:"bitch",5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !      0        array2='{"beauty":2,4:"baker",5:"bitch",5�_�  �  �          �      #    ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !      .        array2='{"beauty":2,"baker",5:"bitch",5�_�  �  �          �      (    ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !      0        array2='{"beauty":2,"baker":4,5:"bitch",5�_�  �  �          �      -    ����                                                                                                                                                                                                                                                                                                                                                V       aD�     �         !      .        array2='{"beauty":2,"baker":4,"bitch",5�_�  �  �          �      5    ����                                                                                                                                                                                                                                                                                                                                                V       aD��     �         !      7                    6:"betray",8:"brazzen",21:"brink"};5�_�  �  �          �      .    ����                                                                                                                                                                                                                                                                                                                                                V       aD��     �         !      :                    6:"betray",8:"brazzen",21:"brink":21};5�_�  �  �          �      !    ����                                                                                                                                                                                                                                                                                                                                                V       aD��     �         !      9                    6:"betray",8:"brazzen":8,"brink":21};5�_�  �  �          �          ����                                                                                                                                                                                                                                                                                                                                                V       aD��     �         !      7                    6:"betray","brazzen":8,"brink":21};5�_�  �              �          ����                                                                                                                                                                                                                                                                                                                                                V       aD��   	 �         !      9                    6:"betray":6,"brazzen":8,"brink":21};5�_�  �          �  �          ����                                                                                                                                                                                                                                                                                                                                                v       aD�     �         "              oreach(array3[i])5�_�  �          �  �           ����                                                                                                                                                                                                                                                                                                                                         
       v       aD�     �         "              $disp5�_�  >          @  ?   (       ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aD��     �   '   )   +      �        <<<<<<<                                                                                                                                                                 string f;5�_�   �           �   �   &   	    ����                                                                                                                                                                                                                                                                                                                                       ,   	       v   	    aDܼ     �   %   '   +      �         <<<<<<<<<<                                                                                                                                                  // last() : Get the last element in the array5�_�      	       
             ����                                                                                                                                                                                                                                                                                                                                       &   	       v   	    aD��     �         $                 }        // size() : Print the number of items in the given dynamic uuuu$display ("fruits_l0.size() = %0d", fruits_l0.size());5�_�                  	          ����                                                                                                                                                                                                                                                                                                                                       %   	       v   	    aD��     �      	   %    5��