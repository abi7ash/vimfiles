Vim�UnDo� s���4Sﰀ���8�T"T����b�414�   )   X        $display("Push_back ahen fruits=%p \n size of fruits=%0d",fruits,fruits.size());   %         x       x   x   x    aP��    _�                             ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �                 class Register;       string name;       rand bit [3:0] rank;       rand bit [3:0] pages;           function new (string name);           this.name=name;       endfunction           function void print();   ?        $display("name=%s rank=%0d pages=%0d",name,rank,pages);       endfunction       endclass    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �                  5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �         $          Register rt[4];   G    string name_arr[4] = '{"alexa","siri","google home","cortana"};               int array[4]='{1,2,3,4};       int res[$];           initial begin5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �                   initial begin5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �                5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �               #//Create a queue to store a strings5�_�      
           	      !    ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �               !//Create a queue to store strings5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �                	//string 5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �                string 5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aP�     �         !      string fruits[$]={"","",""};5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aP�     �         !      "string fruits[$]={"orange","",""};5�_�                       $    ����                                                                                                                                                                                                                                                                                                                                                  v        aP�     �         !      'string fruits[$]={"orange","apple",""};5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aP�$     �         !      ;        $display("----------- Initial Values -----------");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       aP�>     �         !      ;        $display("----------- Initial Values -----------");           foreach(rt[i]) begin   &            rt[i] = new (name_arr[i]);               rt[i].randomize();               rt[i].print();           end       9        $display("----------- Sort by name -----------");   !        rt.sort(x) with (x.name);           foreach(rt[i])                rt[i].print();       @        $display("----------- Sort by rank, pages -----------");   -        rt.sort(x) with ( {x.rank, x.pages});           foreach(rt[i])               rt[i].print();           !        //Array reduction methods   &        $display("array  = %p",array);   +        $display("sum   =%0d",array.sum());        1        $display("prroduct=%0d",array.product());   ,       $display("and   =0x%0h",array.and());   +        $display("or   =0x%0h",array.or());5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       aP�B     �                *        display("or   =0x%0h",array.or());5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       aP�D     �               -        $display("xor   =0x%0h",array.xor());5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       aP�L     �         	              5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       aP�S     �         	              foreach()5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       aP�\     �         	      -        $display("xor   =0x%0h",array.xor());5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       aP�h     �         	      4        $display("fruits[%0d   =0x%0h",array.xor());5�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                v       aP�m     �         	      5        $display("fruits[%0d]   =0x%0h",array.xor());5�_�                       $    ����                                                                                                                                                                                                                                                                                                                                                v       aP�q     �         	      3        $display("fruits[%0d]   =%0h",array.xor());5�_�                       %    ����                                                                                                                                                                                                                                                                                                                                                v       aP�y     �         	      2        $display("fruits[%0d]   =%s",array.xor());5�_�                       2    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �      
   	      2        $display("fruits[%0d]   =%s",i,fruits[i]);5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �      
                 $display()5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �      
                 $display("")5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �      
                 $display("");5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �      
                 $display("fruits=%p");5�_�                     	   %    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �               %        $display("fruits=%p",fruits);5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                       $display()5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                       $display();5�_�   !   #           "          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                       $display("");5�_�   "   $           #      +    ����                                                                                                                                                                                                                                                                                                                                                v       aP��    �               -        $display("Afer deletion, fruits=%p");5�_�   #   %           $      *    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �               ,string fruits[$]={"orange","apple","gauva"};5�_�   $   &           %      C    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �               Jstring fruits[$]={"orange","apple","gauva","kiwi","mango","banana",pear"};5�_�   %   '           &      K    ����                                                                                                                                                                                                                                                                                                                                                v       aP�      �               Kstring fruits[$]={"orange","apple","gauva","kiwi","mango","banana","pear"};5�_�   &   (           '      4    ����                                                                                                                                                                                                                                                                                                                                                v       aP�
     �               4        $display("Afer deletion, fruits=%p",fruits);5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                v       aP�+     �                       $display()5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                v       aP�,     �                       $display("")5�_�   )   +           *      +    ����                                                                                                                                                                                                                                                                                                                                                v       aP�@     �               ,        $display("size of queue fruits=%0d")5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                v       aP�Q     �               /        $display("size of queue fruits=%0d",fr)5�_�   +   -           ,      .    ����                                                                                                                                                                                                                                                                                                                                                v       aP�_     �               /        $display("size of queue fruits=%0d",fr)5�_�   ,   .           -      :    ����                                                                                                                                                                                                                                                                                                                                                v       aP�g     �               :        $display("size of queue fruits=%0d",fruits.size())5�_�   -   /           .          ����                                                                                                                                                                                                                                                                                                                                                v       aP�u     �                       fruits.insert()5�_�   .   0           /          ����                                                                                                                                                                                                                                                                                                                                                v       aP�}     �                       fruits.insert(2,"")5�_�   /   1           0      %    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �               %        fruits.insert(2,"jackfruits")5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                       $display()5�_�   1   3           2      H    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �               H        $display("fruits=%p \n size of fruits=%0d",fruits,fruits.size())5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                       fruits.delete()5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                       fruits.delete(3)5�_�   4   6           5           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �             �             5�_�   5   7           6           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                5�_�   6   8           7           ����                                                                                                                                                                                                                                                                                                                                                v       aP�     �             �             5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                                                v       aP�     �             �             5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                v       aP�     �               I        $display("fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                                                v       aP�/     �               M        $display("Pop fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   :   <           ;      I    ����                                                                                                                                                                                                                                                                                                                                                v       aP�@     �               Y        $display("Pop_front, then fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   ;   >           <      e    ����                                                                                                                                                                                                                                                                                                                                                v       aP�R     �               e        $display("Pop_front, then fruits=%p \n size of fruits=%0d",fruits.pop_front(),fruits.size());5�_�   <   ?   =       >      f    ����                                                                                                                                                                                                                                                                                                                                                v       aP�d     �               f        $display("Pop_front, then fruits=%p \n size of fruits=%0d",fruits.pop_front(),fruits.size());i5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                v       aP�v     �               I        $display("fruits=%p \n size of fruits=%0d",fruits,fruits.size());�             5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                v       aP�{     �               J        $display("$fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   @   B           A      G    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �               W        $display("Pop_back then fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   A   C           B      P    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �               `        $display("Pop_back then fruits=%p \n size of fruits=%0d",fruits.pop_back,fruits.size());5�_�   B   D           C      b    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �               b        $display("Pop_back then fruits=%p \n size of fruits=%0d",fruits.pop_back(),fruits.size());5�_�   C   H           D           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                5�_�   D   I   E       H           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �             �             5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                b        $display("Pop_back then fruits=%p \n size of fruits=%0d",fruits.pop_back(),fruits.size());5�_�   I   K           J          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                `        $display("p_back then fruits=%p \n size of fruits=%0d",fruits.pop_back(),fruits.size());5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �                c        $display("Push_back then fruits=%p \n size of fruits=%0d",fruits.pop_back(),fruits.size());5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         !              5�_�   L   N           M          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         !              fruits.push_back()5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         !              fruits.push_back("")5�_�   N   P           O      "    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         !      "        fruits.push_back("grapes")5�_�   O   Q           P      S    ����                                                                                                                                                                                                                                                                                                                                                v       aP�     �         !      c        $display("Push_back then fruits=%p \n size of fruits=%0d",fruits.pop_back(),fruits.size());5�_�   P   R           Q   !   	    ����                                                                                                                                                                                                                                                                                                                                                v       aP�    �                  	endmodule5�_�   Q   S           R           ����                                                                                                                                                                                                                                                                                                                                                v       aP�9     �         !       5�_�   R   T           S           ����                                                                                                                                                                                                                                                                                                                                                v       aP�:     �         "       5�_�   S   U           T           ����                                                                                                                                                                                                                                                                                                                                                v       aP�O     �         #       5�_�   T   V           U           ����                                                                                                                                                                                                                                                                                                                                                v       aP�Y     �         $       5�_�   U   W           V           ����                                                                                                                                                                                                                                                                                                                                                v       aP�\    �         %       5�_�   V   Y           W          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         %              fruits = fruits2;5�_�   W   Z   X       Y           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         %       5�_�   Y   [           Z           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         &    �         &    5�_�   Z   \           [          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         '              fruits2 = fruits;5�_�   [   ]           \           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         '       5�_�   \   ^           ]           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �   
      (      %        $display("fruits=%p",fruits);   i�         (      i5�_�   ]   _           ^      &    ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �   
      '      &        $display("fruits=%p",fruits);i5�_�   ^   `           _           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         )    �         )    5�_�   _   a           `           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         *       5�_�   `   b           a           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         *      -5�_�   a   c           b           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         *       5�_�   b   d           c           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         *       5�_�   c   e           d           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         *       5�_�   d   f           e           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         *       5�_�   e   g           f           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         *       5�_�   f   h           g           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         )                  fruits={};�         *           �         *       5�_�   g   i           h      *    ����                                                                                                                                                                                                                                                                                                                                                v       aP�     �         (      4        $display("Afer deletion, fruits=%p",fruits);5�_�   h   j           i      @    ����                                                                                                                                                                                                                                                                                                                                                v       aP�     �         (      B        $display("Afer deletion, fruits=%p \n fruits2=%p",fruits);5�_�   i   k           j           ����                                                                                                                                                                                                                                                                                                                                                v       aP�%     �         (    �         (    5�_�   j   l           k          ����                                                                                                                                                                                                                                                                                                                                                v       aP�,    �         )      J        $display("Afer deletion, fruits=%p \n fruits2=%p",fruits,fruits2);5�_�   k   m           l          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         )      I        $display("fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                                                v       aP��    �         )      I        $display("fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   m   p           n           ����                                                                                                                                                                                                                                                                                                                                                v       aP�:     �      !   )      e        $display("Pop_front, then fruits=%p \n size of fruits=%0d",fruits.pop_front(),fruits.size());5�_�   n   q   o       p           ����                                                                                                                                                                                                                                                                                                                                                v       aP�T     �      !   )      h        $display("Pop_front=%p, then fruits=%p \n size of fruits=%0d",fruits.pop_front(),fruits.size());5�_�   p   r           q       Y    ����                                                                                                                                                                                                                                                                                                                                                v       aP�[     �      !   )      h        $display("Pop_front=%p, then fruits=%p \n size of fruits=%0d",fruits.pop_front(),fruits.size());5�_�   q   s           r   "       ����                                                                                                                                                                                                                                                                                                                                                v       aP�m     �   !   #   )      b        $display("Pop_back then fruits=%p \n size of fruits=%0d",fruits.pop_back(),fruits.size());5�_�   r   t           s   "   V    ����                                                                                                                                                                                                                                                                                                                                                v       aP�y    �   !   #   )      e        $display("Pop_back=%p then fruits=%p \n size of fruits=%0d",fruits.pop_back(),fruits.size());5�_�   s   w           t   %       ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �   $   &   )      X        $display("Push_back then fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   t   x   u       w   %       ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �   $   &   )      X        $display("Push_back ahen fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   w               x   %       ����                                                                                                                                                                                                                                                                                                                                                v       aP��    �   $   &   )      X        $display("Push_back then fruits=%p \n size of fruits=%0d",fruits,fruits.size());5�_�   t   v       w   u   %       ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �   %   &   )    �   %   &   )      J        $display("Afer deletion, fruits=%p \n fruits2=%p",fruits,fruits2);5�_�   u               v   &       ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �   %   '   *      I        $displa("Afer deletion, fruits=%p \n fruits2=%p",fruits,fruits2);5�_�   n           p   o           ����                                                                                                                                                                                                                                                                                                                                                v       aP�D     �      !   )      j        $display("Pop_front=%p,\n then fruits=%p \n size of fruits=%0d",fruits.pop_front(),fruits.size());5�_�   W           Y   X           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �         %          	        P5�_�   D   F       H   E           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �             �               $5�_�   E   G           F           ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �             �               $$5�_�   F               G          ����                                                                                                                                                                                                                                                                                                                                                v       aP��     �             �               $$$5�_�   <           >   =          ����                                                                                                                                                                                                                                                                                                                                                v       aP�X     �               e        display("Pop_front, then fruits=%p \n size of fruits=%0d",fruits.pop_front(),fruits.size());i5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �      	        5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �               5��