Vim�UnDo� ���{��	�Y�L�y���"�p�W5be�3�   +           user_st_fruit fruit2;             S       S   S   S    aQZ�    _�                             ����                                                                                                                                                                                                                                                                                                                                                  v        aQ4�     �         0      typedef string str_da [];       class Fruit;       string name;       '    function new(string name="Unkown");           this.name = name;       endfunction   endclass               
module tb;5�_�                            ����                                                                                                                                                                                                                                                                                                                                       #           v        aQ4�     �         $   !   Fruit list[$];       str_da list2[$];   str_da marvel;   str_da dcverse;       initial begin   &        static Fruit f = new("Apple");           list.push_back(f);               f = new("Banana");           list.push_back(f);               foreach(list[i])   8                $display("list[%0d]=%s",i,list[i].name);       !        $display("list=%p",list);           !        //Queue of dynamic arrays   D        marvel = '{"Spiderman","hulk","Captain America","Iron Man"};   5        dcverse = '{"Batman","Wonder Woman","Flash"};                list2.push_back(marvel);   !        list2.push_back(dcverse);               foreach(list2[i])                foreach(list2[i][j])   ?                $display("list2[%0d][%0d]=%s",i,j,list2[i][j]);       %        $display("list2 = %p",list2);               end5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aQ4�     �                   end5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aQ4�     �                 	endmodule5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aQ4�     �                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aQ4�     �                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aQ5     �   
             5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                  v        aQ5"     �                       $display();5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                  v        aQ5$     �                       $display("");5�_�   	              
           ����                                                                                                                                                                                                                                                                                                                                                  v        aQ5,     �               "        $display("st_fruit = %p");5�_�   
                    +    ����                                                                                                                                                                                                                                                                                                                                                  v        aQ51     �               +        $display("st_fruit = %p",st_fruit);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aQ5u     �                       $display()5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aQ5w     �                       $display("")5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aQ5y     �                       $display("");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aQ5�    �                        $display("st_fruit=%p");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aQ5�    �               )        $display("st_fruit=%p",st_fruit);5�_�                    	        ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6     �                5�_�                    
        ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6#     �   	                5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6%     �   	                    �   
          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6*     �   	                struct{5�_�                           ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ61     �                   }st_fruit;5�_�                            ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6S     �                5�_�                            ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6X     �                    �                5�_�                            ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6Z     �                   end5�_�                            ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6]     �                5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6o     �               5        //Adding and using userdefined typedf structs5�_�                       ,    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6p     �               5        //Adding and using userdefined typedf structs5�_�                       6    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6s     �               6        //Adding and using userdefined typedef structs5�_�                           ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �               $        user_st_fruit fruit1 = fruit5�_�                       '    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �               '        user_st_fruit fruit1 = st_fruit5�_�                            ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �         !              $display()5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �         !              $display("")5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �         !              $display("");5�_�   !   #           "      )    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �         !      +        $display("fruit1 = %p\nfruit2=%p");5�_�   "   $           #           ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �      !   !       5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �      "   "              5�_�   $   '           %   !        ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �   !   #   $    �   !   "   $    5�_�   %   (   &       '   "       ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �   !   #   %      9        $display("fruit1 = %p\nfruit2=%p",fruit1,fruit2);5�_�   '   )           (   #        ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ7     �   "   %   %       5�_�   (   *           )   #        ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ7     �   !   #   &      P        $display("puttung fruit1 in fruit2\nit1 = %p\nfruit2=%p",fruit1,fruit2);   i�   "   $   &      i5�_�   )   +           *   "       ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ7     �   !   #   %      R        $display("puttung fruit1 in fruit2\nit1 = %p\nfruit2=%p",fruit1,fruit2);ii5�_�   *   ,           +   "       ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ7     �   !   #   %      S        $displiay("puttung fruit1 in fruit2\nit1 = %p\nfruit2=%p",fruit1,fruit2);ii5�_�   +   -           ,   "   R    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ7     �   !   %   %      R        $display("puttung fruit1 in fruit2\nit1 = %p\nfruit2=%p",fruit1,fruit2);ii5�_�   ,   .           -   "       ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ8G     �   !   #   '      P        $display("puttung fruit1 in fruit2\nit1 = %p\nfruit2=%p",fruit1,fruit2);5�_�   -   /           .   #        ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ8p     �   "   $   '       5�_�   .   0           /   $        ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ8�     �   #   &   '       5�_�   /   1           0   %       ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ8�     �   $   &   (              $display()5�_�   0   2           1   %   "    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ8�     �   $   &   (      "        $display("",fruit1,fruit2)5�_�   1   3           2   %       ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ8�    �   $   &   (      #        $display("",fruit1,fruit2);5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQWg     �         (      #        st_fruit = '{"apple",4,15};5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQWl     �         (      $        st_fruit <= '{"apple",4,15};5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQWr    �         (      (        user_st_fruit fruit1 = st_fruit;5�_�   5   @           6      (    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQW�     �         (      )        user_st_fruit fruit1 <= st_fruit;5�_�   6   A   7       @          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX�     �         (              user_st_fruit fruit1;5�_�   @   B           A          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX�     �         (      !        user_st_fruit fruit1='{};5�_�   A   C           B           ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX�     �         (      %        user_st_fruit fruit1='{"",,};5�_�   B   D           C      '    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX�     �         (      *        user_st_fruit fruit1='{"apple",,};5�_�   C   E           D      )    ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX�    �         (      +        user_st_fruit fruit1='{"apple",4,};5�_�   D   F           E   !        ����                                                                                                                                                                                                                                                                                                                                      	           v       aQY     �      !   '              fruit2 = fruit1;�       !           5�_�   E   G           F          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQYB     �         '      -        user_st_fruit fruit1='{"apple",4,15};5�_�   F   H           G          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQYC     �         '      .        user_st_fruit fruit1 ='{"apple",4,15};5�_�   G   I           H           ����                                                                                                                                                                                                                                                                                                                                      	           v       aQY�     �         '       5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQY�     �         (      /        user_st_fruit fruit1 = '{"apple",4,15};5�_�   I   K           J           ����                                                                                                                                                                                                                                                                                                                                                 v       aQY�     �         (       �         (    5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                                      !           v       aQY�     �         +              user_st_fruit fruit2;5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                                      !           v       aQY�     �         +      ,     user_st_fruit fruit1 = '{"apple",4,15};5�_�   L   O           M          ����                                                                                                                                                                                                                                                                                                                                      !           v       aQY�     �          +      /        user_st_fruit fruit1 = '{"apple",4,15};5�_�   M   P   N       O   %   ,    ����                                                                                                                                                                                                                                                                                                                                      !           v       aQZk     �   $   &   +      P        $display("putting fruit1 in fruit2\nit1 = %p\nfruit2=%p",fruit1,fruit2);5�_�   O   Q           P   $        ����                                                                                                                                                                                                                                                                                                                                      !           v       aQZ�     �   #   %   +       5�_�   P   R           Q   +   	    ����                                                                                                                                                                                                                                                                                                                                      !           v       aQZ�     �   *              	endmodule5�_�   Q   S           R   (       ����                                                                                                                                                                                                                                                                                                                                      !           v       aQZ�    �   '   )   +      7        $display("fruit1=%p\nfruit2=%p",fruit1,fruit2);5�_�   R               S           ����                                                                                                                                                                                                                                                                                                                                      !           v       aQZ�    �      !   +              user_st_fruit fruit2;5�_�   M           O   N           ����                                                                                                                                                                                                                                                                                                                                      !           v       aQY�   
 �      !   +              //user_st_fruit fruit2;5�_�   6   8       @   7           ����                                                                                                                                                                                                                                                                                                                                      	           v       aQW�     �         (           5�_�   7   9           8           ����                                                                                                                                                                                                                                                                                                                                      	           v       aQW�    �         )                  fruit1 = st_fruit;5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQW�     �         *      fruit2;�         *      $        user_st_fruit fruit1,fruit2;5�_�   9   ?           :          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX,    �         )      $        user_st_fruit fruit1,fruit2;5�_�   :       ;       ?          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX�     �         )              fruit1 = st_fruit5�_�   :   <       ?   ;          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQXw     �         )              fruit1 = '{apple";5�_�   ;   >           <          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX�     �         )              fruit1 = '{"apple";5�_�   <       =       >          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX�     �         )      %        fruit1 = '{"apple"er_St_fruit5�_�   <           >   =          ����                                                                                                                                                                                                                                                                                                                                      	           v       aQX�    �         )      "        fruit1 = '{"apple",4,115};5�_�   %           '   &   "       ����                                                                                                                                                                                                                                                                                                                                      	           v       aQ6�     �   "   #   %    �   "   #   %      9        $display("fruit1 = %p\nfruit2=%p",fruit1,fruit2);5��