Vim�UnDo� ���P�ہ�x8IV�M��Z�w�M��\�4��      )        $display("ctrl_reg=%p",ctrl_reg);                             aQ]�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             aQ\"     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �   
                      ctrl_reg = '{};5�_�                       "    ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �   
              "        ctrl_reg = '{4'ha,3'h5,1};5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                         $display()5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                         $display();5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                         $display("");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                          $display("ctrl_reg=%p");5�_�      	                 )    ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                 )        $display("ctrl_reg=%p",ctrl_reg);5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                       ctr;_reg.mode=4'h3;5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                       ctrl_reg.mode=4'h3;5�_�   
                        ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                       $display();5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                       $display("");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                        $display("ctrl_reg=%p");5�_�                       )    ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �               )        $display("ctrl_reg=%p",ctrl_reg);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ\�     �                       $display();5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ]     �                       $display("");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ]     �                        $display("ctrl_reg=%p");5�_�                       )    ����                                                                                                                                                                                                                                                                                                                                                             aQ]     �               )        $display("ctrl_reg=%p",ctrl_reg);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ]    �                   endmodule5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ]q     �               )        $display("ctrl_reg=%p",ctrl_reg);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ]w     �               )        $display("ctrl_reg=%p",ctrl_reg);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             aQ]�     �               )        $display("ctrl_reg=%p",ctrl_reg);5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             aQ]�    �               )        $display("ctrl_reg=%p",ctrl_reg);5��