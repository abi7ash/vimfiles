Vim�UnDo� ț�[���K��S�6G���8�������ʪ��      '            ushorti data=32'hface_cafe;                             aQ�    _�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aQ�     �                  //Create a packed struct   typedef struct packed{       bit [3:0] mode;       bit [2:0] cfg;       bit       en;   	}st_ctrl;       
module tb;       st_ctrl ctrl_reg;       initial begin   "        ctrl_reg = '{4'ha,3'h5,1};   <        $display("Initial contents:\nctrl_reg=%p",ctrl_reg);               ctrl_reg.mode=4'h3;   =        $display("Changing the mode:\nctrl_reg=%p",ctrl_reg);               ctrl_reg=8'hfa;   <        $display("Changing the reg:\nctrl_reg=%p",ctrl_reg);           end       	endmodule    5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aQ�     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aQ�O     �                     typedef enum {};5�_�                       "    ����                                                                                                                                                                                                                                                                                                                                                  v        aQ�U     �                 #    typedef enum {RED,YELLO,GREEN};5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                                  v        aQ�Y     �                 +    typedef enum {RED,YELLO,GREEN} e_light;5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                  v        aQ��     �   
                          $display()5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                  v        aQ��     �   
                          $display("")5�_�   	              
      4    ����                                                                                                                                                                                                                                                                                                                                                  v        aQ��     �   
              5            $display("light=%s\ndata=0x%0h\ncnt=%0d")5�_�   
                    K    ����                                                                                                                                                                                                                                                                                                                                                  v        aQ��     �   
              K            $display("light=%s\ndata=0x%0h\ncnt=%0d",light.name(),data,cnt)5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aQ��     �                       end5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aQ��    �                 	endmodule    �                   end5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aQ�    �               '            ushorti data=32'hface_cafe;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aQ�     �                igned/Create a packed struct5�_�                             ����                                                                                                                                                                                                                                                                                                                                                  v        aQ^c    �                  5��