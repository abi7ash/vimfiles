Vim�UnDo� 3*s�4��e�;C�8_)��gkH�0�6Om�   0   //str_da dcverse;            n       n   n   n    aQ3�    _�                             ����                                                                                                                                                                                                                                                                                                                                                             aP��     �          )      
module tb;5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             aP��     �          *       5�_�                          ����                                                                                                                                                                                                                                                                                                                                       
           v        aP��     �         -          function new()5�_�                       &    ����                                                                                                                                                                                                                                                                                                                                       
           v        aP��     �      	   -      &    function new(string name="Unkown")5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �         1          endfunction5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �         2       5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �   
      2      !//Create a queue to store strings5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �   
             "//Create a queue to storev strings   Kstring fruits[$]={"orange","apple","gauva","kiwi","mango","banana","pear"};       string fruits2[$];    5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �   
      -          initial begin5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �         .      initial begin5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �   
      .          5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP��     �         0           �   
      /          5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP�N     �         /              foreach(fruits[i])5�_�                            ����                                                                                                                                                                                                                                                                                                                                       -           v       aP�b     �                 v        foreach(fruits[i])   2        $display("fruits[%0d]   =%s",i,fruits[i]);       %        $display("fruits=%p",fruits);               fruits2 = fruits;           fruits={};   J        $display("Afer deletion, fruits=%p \n fruits2=%p",fruits,fruits2);               fruits = fruits2;   \        $display("Replicating fruits with fruits2, fruits=%p \n fruits2=%p",fruits,fruits2);               //Queue methods   ;        $display("size of queue fruits=%0d",fruits.size());       &        fruits.insert(2,"jackfruits");   c        $display("After insrtinh jackfruits fruits=%p \n size of fruits=%0d",fruits,fruits.size());                   fruits.delete(3);   l        $display("Deleting element at index 3, now \nfruits=%p \n size of fruits=%0d",fruits,fruits.size());               o        $display("Pop_front=%p, then fruits=%p \n size of fruits=%0d",fruits.pop_front(),fruits,fruits.size());       l        $display("Pop_back=%p then fruits=%p \n size of fruits=%0d",fruits.pop_back(),fruits,fruits.size());       #        fruits.push_back("grapes");   _        $display("Push_back grapes then fruits=%p \n size of fruits=%0d",fruits,fruits.size());        5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aP�k     �                   end5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aP�l     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aP�y     �                       Fruit f = new()5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aP�{     �                       Fruit f = new();5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aP�|    �                       Fruit f = new("");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aQ,�     �                       Fruit f = new("Apple");5�_�      !                      ����                                                                                                                                                                                                                                                                                                                                                  v       aQ,�     �                       list.push_back()5�_�       "           !          ����                                                                                                                                                                                                                                                                                                                                                  v       aQ,�     �                       list.push_back(f)5�_�   !   #           "           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                5�_�   "   $           #           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                �             5�_�   #   %           $           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                Fruit f = new("Apple");5�_�   $   &           %      	    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                         Fruit f = new("Apple");5�_�   %   '           &          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                       Fruit f = new("Apple");5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                       list.push_back(f);5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                       foreach()5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                       foreach(list[i])5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                               $display()5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                               $display();5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ,�     �                               $display("");5�_�   ,   .           -      "    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-     �               %                $display("list[%0d");5�_�   -   /           .      '    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-     �               )                $display("list[%0d]=%s");5�_�   .   0           /      8    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-     �               8                $display("list[%0d]=%s",i,list[i].name);5�_�   /   1           0          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-     �                       $display()5�_�   0   2           1          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-     �                       $display("")5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-#     �                       $display("list=%p")5�_�   2   4           3           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-%    �               !        $display("list=%p",list);    �               !        $display("list=%p",list);    �                        $display("list=%p",list)5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-W    �   
            Fruits list[$];5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-�    �                        Fruit f = new("Banana");5�_�   5   7           6           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ-�     �      
          5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.     �               Fruit list[$];5�_�   7   9           8           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ."     �                   end5�_�   8   :           9           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.#     �                5�_�   9   ;           :           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.&     �                5�_�   :   <           ;      *    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.U     �         !      0        //str_da marvel = '{"Spiderman","hulk","5�_�   ;   =           <      0    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.X     �          !      0        //str_da marvel = '{"Spiderman","hulk","5�_�   <   >           =      
    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.q     �         "      M        //str_da marvel = '{"Spiderman","hulk","Captain America","Iron Man"};5�_�   =   ?           >      
    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.t     �          "              //str5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.v     �          "              str5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �          "      "        str_da dcverse = '{Batman"5�_�   @   B           A      #    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �      "   "      #        str_da dcverse = '{"Batman"5�_�   A   C           B   !       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �       "   $              list2.push_back();5�_�   B   D           C   !        ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �       #   $               list2.push_back(marvel);5�_�   C   E           D   "       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �   !   #   %              list2.push_back()5�_�   D   F           E   "        ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �   !   %   %               list2.push_back(dcverse)5�_�   E   G           F   $       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �   #   %   '              foreach()5�_�   F   H           G   $       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �   #   &   '              foreach(list[i])5�_�   G   I           H   %       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �   $   &   (                  foreach()5�_�   H   J           I   %       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �   $   '   (                  foreach(list[i][j])5�_�   I   K           J   &       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �   %   '   )                      $display()5�_�   J   L           K   &       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ.�     �   %   '   )                      $display("")5�_�   K   M           L   &   ,    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/     �   %   '   )      -                $display("list[%0d][%0d]=%s")5�_�   L   N           M   &   <    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/	     �   %   )   )      <                $display("list[%0d][%0d]=%s",i,j,list[i][j])5�_�   M   O           N   (       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/     �   '   )   +              $display()5�_�   N   P           O   (       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/     �   '   )   +              $display("list = %p)5�_�   O   Q           P   (   "    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/     �   '   *   +      "        $display("list = %p",list)5�_�   P   R           Q   	        ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/R     �      
   ,      typedef string str_da [];5�_�   Q   S           R           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/U     �          ,      class Fruit;5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/W     �          -      i5�_�   S   U           T           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/Z    �         .    �         .    5�_�   T   V           U          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/�     �         /              Fruit f = new("Apple");5�_�   U   W           V          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/�     �         /      $        Fruit tatic  = new("Apple");5�_�   V   X           W          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/�     �         /      %        Fruit static  = new("Apple");5�_�   W   Y           X          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/�     �         /              Fruit  = new("Apple");5�_�   X   Z           Y          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ/�    �         /      %        static Fruit  = new("Apple");5�_�   Y   [           Z   !       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ2�    �       "   /      K        str_da marvel = '{"Spiderman","hulk","Captain America","Iron Man"};5�_�   Z   \           [   !       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ2�     �       "   /      L        str_da marvel <= '{"Spiderman","hulk","Captain America","Iron Man"};5�_�   [   ]           \           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ2�     �         /       5�_�   \   ^           ]   "       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ2�     �   !   #   0      K        str_da marvel = '{"Spiderman","hulk","Captain America","Iron Man"};5�_�   ]   _           ^   #       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ2�   	 �   "   $   0      <        str_da dcverse = '{"Batman","Wonder Woman","Flash"};5�_�   ^   `           _   (       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3     �   '   )   0              foreach(list[i])5�_�   _   a           `   )       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3     �   (   *   0                  foreach(list[i][j])5�_�   `   b           a   *       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3     �   )   +   0      =                $display("list[%0d][%0d]=%s",i,j,list[i][j]);5�_�   a   c           b   *   6    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3     �   )   +   0      >                $display("list2[%0d][%0d]=%s",i,j,list[i][j]);5�_�   b   d           c   ,   !    ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3     �   +   -   0      #        $display("list = %p",list);5�_�   c   e           d   ,       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3   
 �   +   -   0      $        $display("list = %p",list2);5�_�   d   f           e   "       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3M     �   !   #   0      D        marvel = '{"Spiderman","hulk","Captain America","Iron Man"};5�_�   e   g           f   #       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3V     �   "   $   0      5        dcverse = '{"Batman","Wonder Woman","Flash"};5�_�   f   h           g           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3`     �         0      str_da marvel;5�_�   g   i           h           ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3a    �         0      str_da dcverse;5�_�   h   j           i   "       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3�     �   !   #   0      R        static str_da marvel = '{"Spiderman","hulk","Captain America","Iron Man"};5�_�   i   k           j   #       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3�    �   "   $   0      C        static str_da dcverse = '{"Batman","Wonder Woman","Flash"};5�_�   j   l           k   "       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3�     �   !   #   0      K        str_da marvel = '{"Spiderman","hulk","Captain America","Iron Man"};5�_�   k   m           l   #       ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3�     �   "   $   0      <        str_da dcverse = '{"Batman","Wonder Woman","Flash"};5�_�   l   n           m          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3�     �         0      //str_da marvel;5�_�   m               n          ����                                                                                                                                                                                                                                                                                                                                                 v       aQ3�    �         0      //str_da dcverse;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                  v       aP     �           6           Fruit f = new("Apple");                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	        u5�_�      
                    ����                                                                                                                                                                                                                                                                                                                                                             aP��     �         -      %    function new(stringname="Unkown")5�_�                
      $    ����                                                                                                                                                                                                                                                                                                                                       
           v        aP�{     �         -      %    function new(stringname="Unkown"r5�_�   
                    $    ����                                                                                                                                                                                                                                                                                                                                       
           v        aP�|     �         -      %    function new(stringname="Unkown"r5�_�                        $    ����                                                                                                                                                                                                                                                                                                                                       
           v        aP��     �         -      %    function new(stringname="Unkown"u5�_�             
         %    ����                                                                                                                                                                                                                                                                                                                                                             aP��     �         -      &    function new(stringname="Unkown");           this.name=name;       endfunction   endclass        5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             aP�X     �   
      2      !//Create a queue to store strings5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             aP�\     �   
      2       5�_�      	                     ����                                                                                                                                                                                                                                                                                                                                                  v        aP�l     �         2      Kstring fruits[$]={"orange","apple","gauva","kiwi","mango","banana","pear"};5�_�                  	           ����                                                                                                                                                                                                                                                                                                                                                  v        aP�p     �   
      2      Frui5�_�                            ����                                                                                                                                                                                                                                                                                                                                                  v        aP�b     �              5��