Vim�UnDo� ����w�dQ���2�>6Ɨ��f��Nɨ"E��H   9   \        $display("\n\nnow added a new element '6' to id alone.\nid=%p \narray=%p",id,array);   5         �       �   �   �    aD��    _�                            ����                                                                                                                                                                                                                                                                                                                                                            aD�     �                   fruits.5�_�                            ����                                                                                                                                                                                                                                                                                                                                                            aD�     �                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�     �               =    //create a dynamic array that can hold a string of values5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�     �                   fruits=new(3);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�     �   
            +    //create dynamic array to hold 5 values5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�      �                       5�_�      	                      ����                                                                                                                                                                                                                                                                                                                                                            aD�*     �                5�_�      
           	          ����                                                                                                                                                                                                                                                                                                                                                            aD�+     �               i5�_�   	              
          ����                                                                                                                                                                                                                                                                                                                                                            aD�F     �               -        fruits = '{'apple','orange','mango'};5�_�   
                    	    ����                                                                                                                                                                                                                                                                                                                                                            aD�G     �               .        ifruits = '{'apple','orange','mango'};5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�I     �                        5�_�                       -    ����                                                                                                                                                                                                                                                                                                                                                            aD�W     �                -        fruits = '{'apple','orange','mango'};5�_�                       0    ����                                                                                                                                                                                                                                                                                                                                                            aD��     �         #      1        $display("size of fruits is %0d",sizeof()5�_�                       7    ����                                                                                                                                                                                                                                                                                                                                                            aD��     �         #      7        $display("size of fruits is %0d",sizeof(fruits)5�_�                       7    ����                                                                                                                                                                                                                                                                                                                                                            aD��     �         #      8        $display("size of fruits is %0d",sizeof(fruits);5�_�                       9    ����                                                                                                                                                                                                                                                                                                                                                            aD��    �      "   #      9        $display("size of fruits is %0d",sizeof(fruits));5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�D     �         &              fruits=new(3);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�F     �         &              fruits=new[3);5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�K     �         &      -        fruits = '{'apple','orange','mango'};5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�M     �         &      -        fruits = '{"apple','orange','mango'};5�_�                           ����                                                                                                                                                                                                                                                                                                                                                            aD�O     �         &      -        fruits = '{"apple",'orange','mango'};5�_�                       #    ����                                                                                                                                                                                                                                                                                                                                                            aD�R     �         &      -        fruits = '{"apple","orange','mango'};5�_�                       %    ����                                                                                                                                                                                                                                                                                                                                                            aD�S     �         &      -        fruits = '{"apple","orange",'mango'};5�_�                       +    ����                                                                                                                                                                                                                                                                                                                                                            aD�V     �         &      -        fruits = '{"apple","orange","mango'};5�_�                       0    ����                                                                                                                                                                                                                                                                                                                                                            aD�]     �         &      9        $display("size of fruits is %0d",sizeof(fruits));5�_�                       0    ����                                                                                                                                                                                                                                                                                                                                                            aD�c     �         &      2        $display("size of fruits is %0d",fruits));5�_�                    !   *    ����                                                                                                                                                                                                                                                                                                                                                            aD�s     �       %   &      *        $display("\nfruits=%0s\n",fruits);5�_�                    $       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �   #   %   )              fruits.delete();5�_�                    $   #    ����                                                                                                                                                                                                                                                                                                                                                            aD��     �   #   %   )      $        $display("",fruits.delete();5�_�                     $       ����                                                                                                                                                                                                                                                                                                                                                            aD��    �   #   %   )      %        $display("",fruits.delete());5�_�      !               $   7    ����                                                                                                                                                                                                                                                                                                                                                            aD�    �   #   &   (      7        $display("fruits.delete()=%s",fruits.delete());    �   #   %   )      7        $display("fruits.delete()=%s",fruits.delete());    �   #   %   )      7        $display("fruits.delete()=%s",fruits.delete());5�_�       "           !   $       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �   #   &   (      7        $display("fruits.delete()=%s",fruits.delete());5�_�   !   #           "   $       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �   #   %   )              5�_�   "   $           #   %       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �   $   &   )      7        $display("fruits.delete()=%s",fruits.delete());5�_�   #   %           $   %   1    ����                                                                                                                                                                                                                                                                                                                                                            aD��     �   $   &   )      5        $display("fruits.size()=%s",fruits.delete());5�_�   $   &           %   %   "    ����                                                                                                                                                                                                                                                                                                                                                            aD�    �   $   &   )      3        $display("fruits.size()=%s",fruits.size());5�_�   %   '           &   !       ����                                                                                                                                                                                                                                                                                                                                                            aD�z     �       "   )      *        $display("\nfruits=%0s\n",fruits);5�_�   &   (           '   !       ����                                                                                                                                                                                                                                                                                                                                                            aD�|     �       "   )      +        $display("\n fruits=%0s\n",fruits);5�_�   '   )           (   !       ����                                                                                                                                                                                                                                                                                                                                                            aD��    �       "   )      ,        $display("\n fruits=%0s \n",fruits);5�_�   (   *           )   !       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �       "   )      +        $display("\n fruits=%s \n",fruits);5�_�   )   +           *   !       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �       "   )      1        $display("\n ize of ruits=%s \n",fruits);5�_�   *   ,           +   !       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �       "   )      2        $display("\ns ize of ruits=%s \n",fruits);5�_�   +   -           ,   !       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �       "   )      3        $display("\n s ize of ruits=%s \n",fruits);5�_�   ,   .           -   !       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �       "   )      2        $display("\n size of ruits=%s \n",fruits);5�_�   -   /           .   !       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �       "   )      3        $display("\n size of iruits=%s \n",fruits);5�_�   .   0           /   !       ����                                                                                                                                                                                                                                                                                                                                                            aD��     �       "   )      4        $display("\n size of firuits=%s \n",fruits);5�_�   /   1           0   !   &    ����                                                                                                                                                                                                                                                                                                                                                            aD��     �       "   )      3        $display("\n size of fruits=%s \n",fruits);5�_�   0   2           1   !   2    ����                                                                                                                                                                                                                                                                                                                                                            aD��     �       "   )      4        $display("\n size of fruits=%0d \n",fruits);5�_�   1   3           2   !   8    ����                                                                                                                                                                                                                                                                                                                                                            aD��    �       "   )      :        $display("\n size of fruits=%0d \n",fruits.size();5�_�   2   4           3           ����                                                                                                                                                                                                                                                                                                                                                            aD�     �         )       5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                            aD�      �         )              $display();5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                                            aD�#     �         )              $display("");5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                                            aD�4     �         )              $display("fruits[0]");5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                            aD�:     �         )      !        $display("fruits[0]=%s");5�_�   7   9           8      +    ����                                                                                                                                                                                                                                                                                                                                                            aD�?     �         )      +        $display("fruits[0]=%s",fruits[0]);5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                            aD�L     �         *      +        $display("fruits[0]=%s",fruits[0]);5�_�   9   ;           :      $    ����                                                                                                                                                                                                                                                                                                                                                            aD�R     �         *      1        $display("\n \n fruits[0]=%s",fruits[0]);5�_�   :   <           ;   &   !    ����                                                                                                                                                                                                                                                                                                                                                            aD�b    �   %   '   *      3        $display("fruits.size()=%d",fruits.size());5�_�   ;   =           <      !    ����                                                                                                                                                                                                                                                                                                                                                            aD�|     �         *      5        $display("\n \n fruits[0]=%s\n\n",fruits[0]);5�_�   <   >           =      0    ����                                                                                                                                                                                                                                                                                                                                                            aD��    �         *      2        $display("\n \n fruits=%s\n\n",fruits[0]);5�_�   =   ?           >           ����                                                                                                                                                                                                                                                                                                                                                            aD��     �         *      /        $display("\n \n fruits=%s\n\n",fruits);�         *    5�_�   >   @           ?      !    ����                                                                                                                                                                                                                                                                                                                                                            aD��     �         *      0        $display("\n \n fruits=%sf\n\n",fruits);5�_�   ?   A           @      "    ����                                                                                                                                                                                                                                                                                                                                                            aD��   	 �         *      0        $display("\n \n fruits=%pf\n\n",fruits);5�_�   @   B           A   !       ����                                                                                                                                                                                                                                                                                                                           !          #           v       aD��     �       "   *      /        //print the content of the array fruits   ;        $display("\n size of fruits=%0d \n",fruits.size());       *        //delete the contents of the array5�_�   A   C           B   !       ����                                                                                                                                                                                                                                                                                                                           !          !          v       aD��     �       "   '      2                //delete the contents of the array5�_�   B   D           C   #       ����                                                                                                                                                                                                                                                                                                                           !          !          v       aD��     �   "   $   '      4        $display("fruits.size()=%0d",fruits.size());5�_�   C   E           D   #   -    ����                                                                                                                                                                                                                                                                                                                           !          !          v       aD�      �   "   $   '      N        $display("After doing fuits.delete()fruits.size()=%0d",fruits.size());5�_�   D   F           E   #   ,    ����                                                                                                                                                                                                                                                                                                                           !          !          v       aD�   
 �   "   $   '      N        $display("After doing fuits.delete()fruits.size()=%0d",fruits.size());5�_�   E   G           F   #   ?    ����                                                                                                                                                                                                                                                                                                                           !          !          v       aD�     �   "   $   '      P        $display("After doing fuits.delete(), fruits.size()=%0d",fruits.size());5�_�   F   H           G   #       ����                                                                                                                                                                                                                                                                                                                           !          !          v       aD�&    �   "   $   '      T        $display("After doing fuits.delete(), fruits.size()=%0d\n\n",fruits.size());5�_�   G   I           H          ����                                                                                                                                                                                                                                                                                                                           !          !          v       aD�F     �         '      "        //print the array contents5�_�   H   J           I          ����                                                                                                                                                                                                                                                                                                                           !          !          v       aD�J     �         '              //print the contents5�_�   I   K           J          ����                                                                                                                                                                                                                                                                                                                           !          !          v       aD�T     �         '                  array[i]=0;5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                           "          "          v       aD�a     �         (                  $display()5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                           "          "          v       aD�b     �         (                  $display("")5�_�   L   N           M          ����                                                                                                                                                                                                                                                                                                                           "          "          v       aD�h     �         (                   $display("array[%d")5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                           "          "          v       aD�s     �         (      %            $display("array[%d]=%0d")5�_�   N   P           O      %    ����                                                                                                                                                                                                                                                                                                                           "          "          v       aD�v     �         (      &            $display("array[%0d]=%0d")5�_�   O   Q           P      1    ����                                                                                                                                                                                                                                                                                                                           "          "          v       aD�~     �         (      1            $display("array[%0d]=%0d",i,array[i])5�_�   P   R           Q          ����                                                                                                                                                                                                                                                                                                                           "          "          v       aD��     �         (      2            $display("array[%0d]=%0d",i,array[i]);5�_�   Q   S           R      H    ����                                                                                                                                                                                                                                                                                                                           "          "          v       aD��     �         (      H            array[i]=($random%100<0) ?(-1*($random%100)) : $random%100 ;5�_�   R   T           S          ����                                                                                                                                                                                                                                                                                                                           #          #          v       aD��     �         )                  $display();5�_�   S   U           T          ����                                                                                                                                                                                                                                                                                                                           #          #          v       aD��     �         )                  $display("");5�_�   T   V           U      D    ����                                                                                                                                                                                                                                                                                                                           #          #          v       aD��     �         )      J            $display("Adding a random value less than 100 to array[%d]=");5�_�   U   W           V      H    ����                                                                                                                                                                                                                                                                                                                           #          #          v       aD��     �         )      K            $display("Adding a random value less than 100 to array[%0d]=");5�_�   V   X           W      L    ����                                                                                                                                                                                                                                                                                                                           #          #          v       aD��     �         )      N            $display("Adding a random value less than 100 to array[%0d]=%0d");5�_�   W   Y           X      M    ����                                                                                                                                                                                                                                                                                                                           #          #          v       aD��     �         )      R            $display("Adding a random value less than 100 to array[%0d]=%0d",[i]);5�_�   X   Z           Y      M    ����                                                                                                                                                                                                                                                                                                                           #          #          v       aD��     �         )      W            $display("Adding a random value less than 100 to array[%0d]=%0d",array[i]);5�_�   Y   [           Z      M    ����                                                                                                                                                                                                                                                                                                                           #          #          v       aD��    �         )      X            $display("Adding a random value less than 100 to array[%0d]=%0d",,array[i]);5�_�   Z   \           [      %    ����                                                                                                                                                                                                                                                                                                                           #          #          v       aD��     �         )      %        $display("array = %p",array);5�_�   [   ]           \          ����                                                                                                                                                                                                                                                                                                                           $          $          v       aD��     �         *              $display()5�_�   \   ^           ]          ����                                                                                                                                                                                                                                                                                                                           $          $          v       aD��     �         *              $display("")5�_�   ]   _           ^      C    ����                                                                                                                                                                                                                                                                                                                           $          $          v       aD�     �         *      C        $display("Looks like tha value generated is not random...")5�_�   ^   `           _      A    ����                                                                                                                                                                                                                                                                                                                           $          $          v       aD�     �         *      D        $display("Looks like tha value generated is not random...");5�_�   _   a           `      9    ����                                                                                                                                                                                                                                                                                                                           %          %          v       aD�B    �         +      =        it seems to add the same value in each iteration: ");5�_�   `   b           a      V    ����                                                                                                                                                                                                                                                                                                                           %          %          v       aD�W     �         +      Z        it seems to add the same value in each iteration:array = '{-99, 9, 57, 14, 29} ");5�_�   a   c           b      A    ����                                                                                                                                                                                                                                                                                                                           %          %          v       aD�[     �         +      C        $display("Looks like tha value generated is not random...\\5�_�   b   d           c          ����                                                                                                                                                                                                                                                                                                                           %          %          v       aD�^    �         +      E        $display("Looks like tha value generated is not random...\n\\5�_�   c   e           d      G    ����                                                                                                                                                                                                                                                                                                                           %          %          v       aD�r    �         +      E        $display("\nLooks like tha value generated is not random...\n   \        it seems to add the same value in each iteration:array = '{-99, 9, 57, 14, 29}\n ");�         +      G        $display("\nLooks like tha value generated is not random...\n\\5�_�   d   f           e      u    ����                                                                                                                                                                                                                                                                                                                           $          $          v       aD��     �         *      �        $display("\nLooks like tha value generated is not random...\nit seems to add the same value in each iteration:array = '{-99, 9, 57, 14, 29}\n ");5�_�   e   g           f          ����                                                                                                                                                                                                                                                                                                                           $          $          v       aD�4     �         *          int array[];5�_�   f   h           g           ����                                                                                                                                                                                                                                                                                                                           $          $          v       aD�>     �         *       5�_�   g   i           h   )        ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�g     �   (   +   ,       5�_�   h   j           i   )        ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�i     �   (   /   -       5�_�   i   k           j   .       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   -   /   2              $display();5�_�   j   l           k   .       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   -   /   2              $display("");5�_�   k   m           l   .   *    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   -   /   2      ,        $display("id=%p and size of id=%d");5�_�   l   n           m   .   9    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   -   1   2      9        $display("id=%p and size of id=%d",id,id.size());5�_�   m   o           n   0   &    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   /   1   4      2        //increase the size of id and add another 5�_�   n   p           o   0       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   /   2   4              //add another 5�_�   o   q           p   1       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�)     �   0   2   5              id = new[id.size()+1]()5�_�   p   r           q   1   !    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�*     �   0   5   5      !        id = new[id.size()+1](id)5�_�   q   s           r   4       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�X     �   3   5   8               //lets see its contents 5�_�   r   t           s   4       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�`     �   3   5   8              //compare contents 5�_�   s   u           t   4       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�b     �   3   5   8      #        //compare contentsof id an 5�_�   t   v           u   4   $    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�e     �   3   6   8      $        //compare contents of id an 5�_�   u   w           v   5       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�q     �   4   6   9              $display()5�_�   v   x           w   5       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�r     �   4   6   9              $display();5�_�   w   y           x   5       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�t    �   4   6   9              $display("");5�_�   x   z           y   5   $    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��    �   4   6   9      &        $display("id=%p \n array=%p");5�_�   y   {           z   .       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   -   /   9      9        $display("id=%p and size of id=%d",id,id.size());5�_�   z   |           {   .   9    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   -   /   9      `        $display("array contents have been replicated to id=%p and size of id=%d",id,id.size());5�_�   {   }           |   .       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   -   /   9      h        $display("array contents have been replicated to id./nso id=%p and size of id=%d",id,id.size());5�_�   |   ~           }   .   A    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   -   /   9      l        $display("\n\narray contents have been replicated to id./nso id=%p and size of id=%d",id,id.size());5�_�   }              ~   .   [    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   -   /   9      l        $display("\n\narray contents have been replicated to id.\nso id=%p and size of id=%d",id,id.size());5�_�   ~   �              5       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��     �   4   6   9      /        $display("id=%p \n array=%p",id,array);5�_�      �           �   5   5    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�     �   4   6   9      T        $display("now added a new element to id alone\nid=%p \n array=%p",id,array);5�_�   �   �           �   5   *    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�    �   4   6   9      U        $display("now added a new element to id alone.\nid=%p \n array=%p",id,array);5�_�   �   �           �   5   E    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�5     �   4   6   9      Y        $display("now added a new element '6' to id alone.\nid=%p \n array=%p",id,array);5�_�   �   �           �   5       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�;     �   4   6   9      X        $display("now added a new element '6' to id alone.\nid=%p \narray=%p",id,array);5�_�   �   �           �   .   B    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�K     �   -   /   9      m        $display("\n\narray contents have been replicated to id.\nso id=%p and size of id=%0d",id,id.size());5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�Q    �   -   /   9      o        $display("\n\narray contents have been replicated to id.\n\nso id=%p and size of id=%0d",id,id.size());5�_�   �   �           �   .       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�q     �   -   /   9      q        $display("\n\n\narray contents have been replicated to id.\n\nso id=%p and size of id=%0d",id,id.size());5�_�   �   �           �   .   @    ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD�x     �   -   /   9      m        $display("\narray contents have been replicated to id.\n\nso id=%p and size of id=%0d",id,id.size());5�_�   �               �   5       ����                                                                                                                                                                                                                                                                                                                           &          &          v       aD��    �   4   6   9      \        $display("\n\nnow added a new element '6' to id alone.\nid=%p \narray=%p",id,array);5��